--------------------------------------------------------------------------------
--     This file is owned and controlled by Xilinx and must be used           --
--     solely for design, simulation, implementation and creation of          --
--     design files limited to Xilinx devices or technologies. Use            --
--     with non-Xilinx devices or technologies is expressly prohibited        --
--     and immediately terminates your license.                               --
--                                                                            --
--     XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS"          --
--     SOLELY FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR                --
--     XILINX DEVICES.  BY PROVIDING THIS DESIGN, CODE, OR INFORMATION        --
--     AS ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE, APPLICATION            --
--     OR STANDARD, XILINX IS MAKING NO REPRESENTATION THAT THIS              --
--     IMPLEMENTATION IS FREE FROM ANY CLAIMS OF INFRINGEMENT,                --
--     AND YOU ARE RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY REQUIRE       --
--     FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY DISCLAIMS ANY               --
--     WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE                --
--     IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR         --
--     REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF        --
--     INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS        --
--     FOR A PARTICULAR PURPOSE.                                              --
--                                                                            --
--     Xilinx products are not intended for use in life support               --
--     appliances, devices, or systems. Use in such applications are          --
--     expressly prohibited.                                                  --
--                                                                            --
--     (c) Copyright 1995-2004 Xilinx, Inc.                                   --
--     All rights reserved.                                                   --
--------------------------------------------------------------------------------

-- synopsys translate_off
LIBRARY std, ieee;
USE std.standard.ALL;
USE ieee.std_logic_1164.ALL;

LIBRARY unisim;
USE unisim.vcomponents.ALL;


LIBRARY XilinxCoreLib;
USE XilinxCoreLib.c_addsub_v5_0_comp.ALL;
USE XilinxCoreLib.c_da_fir_v7_0_comp.ALL;
USE XilinxCoreLib.c_mux_bus_v5_0_comp.ALL;
USE XilinxCoreLib.c_counter_binary_v5_0_comp.ALL;
USE XilinxCoreLib.c_cic_v3_0_comp.ALL;
USE XilinxCoreLib.c_reg_fd_v5_0_comp.ALL;
USE XilinxCoreLib.c_dds_v4_1_comp.ALL;
USE XilinxCoreLib.c_shift_ram_v5_0_comp.ALL;
USE XilinxCoreLib.mult_gen_v5_0_comp.ALL;
USE XilinxCoreLib.c_gate_bit_v5_0_comp.ALL;

ENTITY ddcv_orig IS
   PORT (
      DIN : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
      ND : IN STD_LOGIC;
      CLK : IN STD_LOGIC;
      ADDR : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      LD_DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      WE : IN STD_LOGIC;
      SEL : IN STD_LOGIC;
      RDY : OUT STD_LOGIC;
      RFD : OUT STD_LOGIC;
      DOUT_I : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
      DOUT_Q : OUT STD_LOGIC_VECTOR(29 DOWNTO 0)   
);
END ddcv_orig;

ARCHITECTURE xilinx OF ddcv_orig IS 

-- Signals for connecting to instantiations
   SIGNAL BU4_I0 : STD_LOGIC;
   SIGNAL BU4_I1 : STD_LOGIC;
   SIGNAL BU4_I2 : STD_LOGIC;
   SIGNAL BU4_I3 : STD_LOGIC;
   SIGNAL BU4_O : STD_LOGIC;
   SIGNAL BU8_I0 : STD_LOGIC;
   SIGNAL BU8_I1 : STD_LOGIC;
   SIGNAL BU8_I2 : STD_LOGIC;
   SIGNAL BU8_I3 : STD_LOGIC;
   SIGNAL BU8_O : STD_LOGIC;
   SIGNAL BU10_I0 : STD_LOGIC;
   SIGNAL BU10_I1 : STD_LOGIC;
   SIGNAL BU10_I2 : STD_LOGIC;
   SIGNAL BU10_I3 : STD_LOGIC;
   SIGNAL BU10_O : STD_LOGIC;
   SIGNAL BU1292_D : STD_LOGIC;
   SIGNAL BU1292_C : STD_LOGIC;
   SIGNAL BU1292_CE : STD_LOGIC;
   SIGNAL BU1292_Q : STD_LOGIC;
   SIGNAL BU14_D : STD_LOGIC;
   SIGNAL BU14_CE : STD_LOGIC;
   SIGNAL BU14_CLK : STD_LOGIC;
   SIGNAL BU14_A0 : STD_LOGIC;
   SIGNAL BU14_A1 : STD_LOGIC;
   SIGNAL BU14_A2 : STD_LOGIC;
   SIGNAL BU14_A3 : STD_LOGIC;
   SIGNAL BU14_Q : STD_LOGIC;
   SIGNAL BU16_D : STD_LOGIC;
   SIGNAL BU16_C : STD_LOGIC;
   SIGNAL BU16_CE : STD_LOGIC;
   SIGNAL BU16_Q : STD_LOGIC;
   SIGNAL BU17_D : STD_LOGIC;
   SIGNAL BU17_CE : STD_LOGIC;
   SIGNAL BU17_CLK : STD_LOGIC;
   SIGNAL BU17_A0 : STD_LOGIC;
   SIGNAL BU17_A1 : STD_LOGIC;
   SIGNAL BU17_A2 : STD_LOGIC;
   SIGNAL BU17_A3 : STD_LOGIC;
   SIGNAL BU17_Q : STD_LOGIC;
   SIGNAL BU19_D : STD_LOGIC;
   SIGNAL BU19_C : STD_LOGIC;
   SIGNAL BU19_CE : STD_LOGIC;
   SIGNAL BU19_Q : STD_LOGIC;
   SIGNAL BU20_D : STD_LOGIC;
   SIGNAL BU20_CE : STD_LOGIC;
   SIGNAL BU20_CLK : STD_LOGIC;
   SIGNAL BU20_A0 : STD_LOGIC;
   SIGNAL BU20_A1 : STD_LOGIC;
   SIGNAL BU20_A2 : STD_LOGIC;
   SIGNAL BU20_A3 : STD_LOGIC;
   SIGNAL BU20_Q : STD_LOGIC;
   SIGNAL BU22_D : STD_LOGIC;
   SIGNAL BU22_C : STD_LOGIC;
   SIGNAL BU22_CE : STD_LOGIC;
   SIGNAL BU22_Q : STD_LOGIC;
   SIGNAL BU23_D : STD_LOGIC;
   SIGNAL BU23_CE : STD_LOGIC;
   SIGNAL BU23_CLK : STD_LOGIC;
   SIGNAL BU23_A0 : STD_LOGIC;
   SIGNAL BU23_A1 : STD_LOGIC;
   SIGNAL BU23_A2 : STD_LOGIC;
   SIGNAL BU23_A3 : STD_LOGIC;
   SIGNAL BU23_Q : STD_LOGIC;
   SIGNAL BU25_D : STD_LOGIC;
   SIGNAL BU25_C : STD_LOGIC;
   SIGNAL BU25_CE : STD_LOGIC;
   SIGNAL BU25_Q : STD_LOGIC;
   SIGNAL BU26_D : STD_LOGIC;
   SIGNAL BU26_CE : STD_LOGIC;
   SIGNAL BU26_CLK : STD_LOGIC;
   SIGNAL BU26_A0 : STD_LOGIC;
   SIGNAL BU26_A1 : STD_LOGIC;
   SIGNAL BU26_A2 : STD_LOGIC;
   SIGNAL BU26_A3 : STD_LOGIC;
   SIGNAL BU26_Q : STD_LOGIC;
   SIGNAL BU28_D : STD_LOGIC;
   SIGNAL BU28_C : STD_LOGIC;
   SIGNAL BU28_CE : STD_LOGIC;
   SIGNAL BU28_Q : STD_LOGIC;
   SIGNAL BU29_D : STD_LOGIC;
   SIGNAL BU29_CE : STD_LOGIC;
   SIGNAL BU29_CLK : STD_LOGIC;
   SIGNAL BU29_A0 : STD_LOGIC;
   SIGNAL BU29_A1 : STD_LOGIC;
   SIGNAL BU29_A2 : STD_LOGIC;
   SIGNAL BU29_A3 : STD_LOGIC;
   SIGNAL BU29_Q : STD_LOGIC;
   SIGNAL BU31_D : STD_LOGIC;
   SIGNAL BU31_C : STD_LOGIC;
   SIGNAL BU31_CE : STD_LOGIC;
   SIGNAL BU31_Q : STD_LOGIC;
   SIGNAL BU32_D : STD_LOGIC;
   SIGNAL BU32_CE : STD_LOGIC;
   SIGNAL BU32_CLK : STD_LOGIC;
   SIGNAL BU32_A0 : STD_LOGIC;
   SIGNAL BU32_A1 : STD_LOGIC;
   SIGNAL BU32_A2 : STD_LOGIC;
   SIGNAL BU32_A3 : STD_LOGIC;
   SIGNAL BU32_Q : STD_LOGIC;
   SIGNAL BU34_D : STD_LOGIC;
   SIGNAL BU34_C : STD_LOGIC;
   SIGNAL BU34_CE : STD_LOGIC;
   SIGNAL BU34_Q : STD_LOGIC;
   SIGNAL BU35_D : STD_LOGIC;
   SIGNAL BU35_CE : STD_LOGIC;
   SIGNAL BU35_CLK : STD_LOGIC;
   SIGNAL BU35_A0 : STD_LOGIC;
   SIGNAL BU35_A1 : STD_LOGIC;
   SIGNAL BU35_A2 : STD_LOGIC;
   SIGNAL BU35_A3 : STD_LOGIC;
   SIGNAL BU35_Q : STD_LOGIC;
   SIGNAL BU37_D : STD_LOGIC;
   SIGNAL BU37_C : STD_LOGIC;
   SIGNAL BU37_CE : STD_LOGIC;
   SIGNAL BU37_Q : STD_LOGIC;
   SIGNAL BU38_D : STD_LOGIC;
   SIGNAL BU38_CE : STD_LOGIC;
   SIGNAL BU38_CLK : STD_LOGIC;
   SIGNAL BU38_A0 : STD_LOGIC;
   SIGNAL BU38_A1 : STD_LOGIC;
   SIGNAL BU38_A2 : STD_LOGIC;
   SIGNAL BU38_A3 : STD_LOGIC;
   SIGNAL BU38_Q : STD_LOGIC;
   SIGNAL BU40_D : STD_LOGIC;
   SIGNAL BU40_C : STD_LOGIC;
   SIGNAL BU40_CE : STD_LOGIC;
   SIGNAL BU40_Q : STD_LOGIC;
   SIGNAL BU41_D : STD_LOGIC;
   SIGNAL BU41_CE : STD_LOGIC;
   SIGNAL BU41_CLK : STD_LOGIC;
   SIGNAL BU41_A0 : STD_LOGIC;
   SIGNAL BU41_A1 : STD_LOGIC;
   SIGNAL BU41_A2 : STD_LOGIC;
   SIGNAL BU41_A3 : STD_LOGIC;
   SIGNAL BU41_Q : STD_LOGIC;
   SIGNAL BU43_D : STD_LOGIC;
   SIGNAL BU43_C : STD_LOGIC;
   SIGNAL BU43_CE : STD_LOGIC;
   SIGNAL BU43_Q : STD_LOGIC;
   SIGNAL BU44_D : STD_LOGIC;
   SIGNAL BU44_CE : STD_LOGIC;
   SIGNAL BU44_CLK : STD_LOGIC;
   SIGNAL BU44_A0 : STD_LOGIC;
   SIGNAL BU44_A1 : STD_LOGIC;
   SIGNAL BU44_A2 : STD_LOGIC;
   SIGNAL BU44_A3 : STD_LOGIC;
   SIGNAL BU44_Q : STD_LOGIC;
   SIGNAL BU46_D : STD_LOGIC;
   SIGNAL BU46_C : STD_LOGIC;
   SIGNAL BU46_CE : STD_LOGIC;
   SIGNAL BU46_Q : STD_LOGIC;
   SIGNAL BU47_D : STD_LOGIC;
   SIGNAL BU47_CE : STD_LOGIC;
   SIGNAL BU47_CLK : STD_LOGIC;
   SIGNAL BU47_A0 : STD_LOGIC;
   SIGNAL BU47_A1 : STD_LOGIC;
   SIGNAL BU47_A2 : STD_LOGIC;
   SIGNAL BU47_A3 : STD_LOGIC;
   SIGNAL BU47_Q : STD_LOGIC;
   SIGNAL BU49_D : STD_LOGIC;
   SIGNAL BU49_C : STD_LOGIC;
   SIGNAL BU49_CE : STD_LOGIC;
   SIGNAL BU49_Q : STD_LOGIC;
   SIGNAL BU50_D : STD_LOGIC;
   SIGNAL BU50_CE : STD_LOGIC;
   SIGNAL BU50_CLK : STD_LOGIC;
   SIGNAL BU50_A0 : STD_LOGIC;
   SIGNAL BU50_A1 : STD_LOGIC;
   SIGNAL BU50_A2 : STD_LOGIC;
   SIGNAL BU50_A3 : STD_LOGIC;
   SIGNAL BU50_Q : STD_LOGIC;
   SIGNAL BU52_D : STD_LOGIC;
   SIGNAL BU52_C : STD_LOGIC;
   SIGNAL BU52_CE : STD_LOGIC;
   SIGNAL BU52_Q : STD_LOGIC;
   SIGNAL BU53_D : STD_LOGIC;
   SIGNAL BU53_CE : STD_LOGIC;
   SIGNAL BU53_CLK : STD_LOGIC;
   SIGNAL BU53_A0 : STD_LOGIC;
   SIGNAL BU53_A1 : STD_LOGIC;
   SIGNAL BU53_A2 : STD_LOGIC;
   SIGNAL BU53_A3 : STD_LOGIC;
   SIGNAL BU53_Q : STD_LOGIC;
   SIGNAL BU55_D : STD_LOGIC;
   SIGNAL BU55_C : STD_LOGIC;
   SIGNAL BU55_CE : STD_LOGIC;
   SIGNAL BU55_Q : STD_LOGIC;
   SIGNAL BU57_DATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
   SIGNAL BU57_WE : STD_LOGIC;
   SIGNAL BU57_CLK : STD_LOGIC;
   SIGNAL BU57_CE : STD_LOGIC;
   SIGNAL BU57_RDY : STD_LOGIC;
   SIGNAL BU57_SINE : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU57_COSINE : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1294_I0 : STD_LOGIC;
   SIGNAL BU1294_I1 : STD_LOGIC;
   SIGNAL BU1294_I2 : STD_LOGIC;
   SIGNAL BU1294_I3 : STD_LOGIC;
   SIGNAL BU1294_O : STD_LOGIC;
   SIGNAL BU1296_clk : STD_LOGIC;
   SIGNAL BU1296_a : STD_LOGIC_VECTOR(13 DOWNTO 0);
   SIGNAL BU1296_b : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1296_o : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1296_q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1296_a_signed : STD_LOGIC;
   SIGNAL BU1296_loadb : STD_LOGIC;
   SIGNAL BU1296_load_done : STD_LOGIC;
   SIGNAL BU1296_swapb : STD_LOGIC;
   SIGNAL BU1296_ce : STD_LOGIC;
   SIGNAL BU1296_aclr : STD_LOGIC;
   SIGNAL BU1296_sclr : STD_LOGIC;
   SIGNAL BU1296_rfd : STD_LOGIC;
   SIGNAL BU1296_nd : STD_LOGIC;
   SIGNAL BU1296_rdy : STD_LOGIC;
   SIGNAL BU1517_I : STD_LOGIC_VECTOR(4 DOWNTO 0);
   SIGNAL BU1517_O : STD_LOGIC;
   SIGNAL BU1526_I0 : STD_LOGIC;
   SIGNAL BU1526_I1 : STD_LOGIC;
   SIGNAL BU1526_I2 : STD_LOGIC;
   SIGNAL BU1526_I3 : STD_LOGIC;
   SIGNAL BU1526_O : STD_LOGIC;
   SIGNAL BU1527_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU1527_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1527_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU1628_I0 : STD_LOGIC;
   SIGNAL BU1628_I1 : STD_LOGIC;
   SIGNAL BU1628_I2 : STD_LOGIC;
   SIGNAL BU1628_I3 : STD_LOGIC;
   SIGNAL BU1628_O : STD_LOGIC;
   SIGNAL BU1630_I0 : STD_LOGIC;
   SIGNAL BU1630_I1 : STD_LOGIC;
   SIGNAL BU1630_I2 : STD_LOGIC;
   SIGNAL BU1630_I3 : STD_LOGIC;
   SIGNAL BU1630_O : STD_LOGIC;
   SIGNAL BU1631_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU1631_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU1631_CLK : STD_LOGIC;
   SIGNAL BU1631_SCLR : STD_LOGIC;
   SIGNAL BU1631_SSET : STD_LOGIC;
   SIGNAL BU1724_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1724_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1724_CLK : STD_LOGIC;
   SIGNAL BU1724_SCLR : STD_LOGIC;
   SIGNAL BU1724_SSET : STD_LOGIC;
   SIGNAL BU1729_CLK : STD_LOGIC;
   SIGNAL BU1729_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1729_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1734_clk : STD_LOGIC;
   SIGNAL BU1734_a : STD_LOGIC_VECTOR(13 DOWNTO 0);
   SIGNAL BU1734_b : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1734_o : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1734_q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1734_a_signed : STD_LOGIC;
   SIGNAL BU1734_loadb : STD_LOGIC;
   SIGNAL BU1734_load_done : STD_LOGIC;
   SIGNAL BU1734_swapb : STD_LOGIC;
   SIGNAL BU1734_ce : STD_LOGIC;
   SIGNAL BU1734_aclr : STD_LOGIC;
   SIGNAL BU1734_sclr : STD_LOGIC;
   SIGNAL BU1734_rfd : STD_LOGIC;
   SIGNAL BU1734_nd : STD_LOGIC;
   SIGNAL BU1734_rdy : STD_LOGIC;
   SIGNAL BU1955_I : STD_LOGIC_VECTOR(4 DOWNTO 0);
   SIGNAL BU1955_O : STD_LOGIC;
   SIGNAL BU1964_I0 : STD_LOGIC;
   SIGNAL BU1964_I1 : STD_LOGIC;
   SIGNAL BU1964_I2 : STD_LOGIC;
   SIGNAL BU1964_I3 : STD_LOGIC;
   SIGNAL BU1964_O : STD_LOGIC;
   SIGNAL BU1965_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU1965_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1965_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU2066_I0 : STD_LOGIC;
   SIGNAL BU2066_I1 : STD_LOGIC;
   SIGNAL BU2066_I2 : STD_LOGIC;
   SIGNAL BU2066_I3 : STD_LOGIC;
   SIGNAL BU2066_O : STD_LOGIC;
   SIGNAL BU2068_I0 : STD_LOGIC;
   SIGNAL BU2068_I1 : STD_LOGIC;
   SIGNAL BU2068_I2 : STD_LOGIC;
   SIGNAL BU2068_I3 : STD_LOGIC;
   SIGNAL BU2068_O : STD_LOGIC;
   SIGNAL BU2069_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2069_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2069_CLK : STD_LOGIC;
   SIGNAL BU2069_SCLR : STD_LOGIC;
   SIGNAL BU2069_SSET : STD_LOGIC;
   SIGNAL BU2162_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2162_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2162_CLK : STD_LOGIC;
   SIGNAL BU2162_SCLR : STD_LOGIC;
   SIGNAL BU2162_SSET : STD_LOGIC;
   SIGNAL BU2457_D : STD_LOGIC;
   SIGNAL BU2457_C : STD_LOGIC;
   SIGNAL BU2457_CE : STD_LOGIC;
   SIGNAL BU2457_Q : STD_LOGIC;
   SIGNAL BU2461_I : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2461_O : STD_LOGIC;
   SIGNAL BU2489_I0 : STD_LOGIC;
   SIGNAL BU2489_I1 : STD_LOGIC;
   SIGNAL BU2489_I2 : STD_LOGIC;
   SIGNAL BU2489_I3 : STD_LOGIC;
   SIGNAL BU2489_O : STD_LOGIC;
   SIGNAL BU2490_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2490_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2490_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU2591_I0 : STD_LOGIC;
   SIGNAL BU2591_I1 : STD_LOGIC;
   SIGNAL BU2591_I2 : STD_LOGIC;
   SIGNAL BU2591_I3 : STD_LOGIC;
   SIGNAL BU2591_O : STD_LOGIC;
   SIGNAL BU2593_I0 : STD_LOGIC;
   SIGNAL BU2593_I1 : STD_LOGIC;
   SIGNAL BU2593_I2 : STD_LOGIC;
   SIGNAL BU2593_I3 : STD_LOGIC;
   SIGNAL BU2593_O : STD_LOGIC;
   SIGNAL BU2594_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2594_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2594_CLK : STD_LOGIC;
   SIGNAL BU2594_SCLR : STD_LOGIC;
   SIGNAL BU2594_SSET : STD_LOGIC;
   SIGNAL BU2687_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2687_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2687_CLK : STD_LOGIC;
   SIGNAL BU2687_SCLR : STD_LOGIC;
   SIGNAL BU2687_SSET : STD_LOGIC;
   SIGNAL BU7487_I : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU7487_O : STD_LOGIC;
   SIGNAL BU7515_I0 : STD_LOGIC;
   SIGNAL BU7515_I1 : STD_LOGIC;
   SIGNAL BU7515_I2 : STD_LOGIC;
   SIGNAL BU7515_I3 : STD_LOGIC;
   SIGNAL BU7515_O : STD_LOGIC;
   SIGNAL BU7516_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU7516_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU7516_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU7617_I0 : STD_LOGIC;
   SIGNAL BU7617_I1 : STD_LOGIC;
   SIGNAL BU7617_I2 : STD_LOGIC;
   SIGNAL BU7617_I3 : STD_LOGIC;
   SIGNAL BU7617_O : STD_LOGIC;
   SIGNAL BU7619_I0 : STD_LOGIC;
   SIGNAL BU7619_I1 : STD_LOGIC;
   SIGNAL BU7619_I2 : STD_LOGIC;
   SIGNAL BU7619_I3 : STD_LOGIC;
   SIGNAL BU7619_O : STD_LOGIC;
   SIGNAL BU7620_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU7620_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU7620_CLK : STD_LOGIC;
   SIGNAL BU7620_SCLR : STD_LOGIC;
   SIGNAL BU7620_SSET : STD_LOGIC;
   SIGNAL BU7713_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU7713_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU7713_CLK : STD_LOGIC;
   SIGNAL BU7713_SCLR : STD_LOGIC;
   SIGNAL BU7713_SSET : STD_LOGIC;
   SIGNAL BU2173_D : STD_LOGIC;
   SIGNAL BU2173_C : STD_LOGIC;
   SIGNAL BU2173_CE : STD_LOGIC;
   SIGNAL BU2173_Q : STD_LOGIC;
   SIGNAL BU2175_D : STD_LOGIC;
   SIGNAL BU2175_C : STD_LOGIC;
   SIGNAL BU2175_CE : STD_LOGIC;
   SIGNAL BU2175_Q : STD_LOGIC;
   SIGNAL BU2177_D : STD_LOGIC;
   SIGNAL BU2177_C : STD_LOGIC;
   SIGNAL BU2177_CE : STD_LOGIC;
   SIGNAL BU2177_Q : STD_LOGIC;
   SIGNAL BU2179_D : STD_LOGIC;
   SIGNAL BU2179_C : STD_LOGIC;
   SIGNAL BU2179_CE : STD_LOGIC;
   SIGNAL BU2179_Q : STD_LOGIC;
   SIGNAL BU2181_D : STD_LOGIC;
   SIGNAL BU2181_C : STD_LOGIC;
   SIGNAL BU2181_CE : STD_LOGIC;
   SIGNAL BU2181_Q : STD_LOGIC;
   SIGNAL BU2183_D : STD_LOGIC;
   SIGNAL BU2183_C : STD_LOGIC;
   SIGNAL BU2183_CE : STD_LOGIC;
   SIGNAL BU2183_Q : STD_LOGIC;
   SIGNAL BU2185_D : STD_LOGIC;
   SIGNAL BU2185_C : STD_LOGIC;
   SIGNAL BU2185_CE : STD_LOGIC;
   SIGNAL BU2185_Q : STD_LOGIC;
   SIGNAL BU2187_D : STD_LOGIC;
   SIGNAL BU2187_C : STD_LOGIC;
   SIGNAL BU2187_CE : STD_LOGIC;
   SIGNAL BU2187_Q : STD_LOGIC;
   SIGNAL BU2189_D : STD_LOGIC;
   SIGNAL BU2189_C : STD_LOGIC;
   SIGNAL BU2189_CE : STD_LOGIC;
   SIGNAL BU2189_Q : STD_LOGIC;
   SIGNAL BU2191_D : STD_LOGIC;
   SIGNAL BU2191_C : STD_LOGIC;
   SIGNAL BU2191_CE : STD_LOGIC;
   SIGNAL BU2191_Q : STD_LOGIC;
   SIGNAL BU2193_D : STD_LOGIC;
   SIGNAL BU2193_C : STD_LOGIC;
   SIGNAL BU2193_CE : STD_LOGIC;
   SIGNAL BU2193_Q : STD_LOGIC;
   SIGNAL BU2195_D : STD_LOGIC;
   SIGNAL BU2195_C : STD_LOGIC;
   SIGNAL BU2195_CE : STD_LOGIC;
   SIGNAL BU2195_Q : STD_LOGIC;
   SIGNAL BU2197_D : STD_LOGIC;
   SIGNAL BU2197_C : STD_LOGIC;
   SIGNAL BU2197_CE : STD_LOGIC;
   SIGNAL BU2197_Q : STD_LOGIC;
   SIGNAL BU2199_D : STD_LOGIC;
   SIGNAL BU2199_C : STD_LOGIC;
   SIGNAL BU2199_CE : STD_LOGIC;
   SIGNAL BU2199_Q : STD_LOGIC;
   SIGNAL BU2201_D : STD_LOGIC;
   SIGNAL BU2201_C : STD_LOGIC;
   SIGNAL BU2201_CE : STD_LOGIC;
   SIGNAL BU2201_Q : STD_LOGIC;
   SIGNAL BU2203_D : STD_LOGIC;
   SIGNAL BU2203_C : STD_LOGIC;
   SIGNAL BU2203_CE : STD_LOGIC;
   SIGNAL BU2203_Q : STD_LOGIC;
   SIGNAL BU2205_D : STD_LOGIC;
   SIGNAL BU2205_C : STD_LOGIC;
   SIGNAL BU2205_CE : STD_LOGIC;
   SIGNAL BU2205_Q : STD_LOGIC;
   SIGNAL BU2207_D : STD_LOGIC;
   SIGNAL BU2207_C : STD_LOGIC;
   SIGNAL BU2207_CE : STD_LOGIC;
   SIGNAL BU2207_Q : STD_LOGIC;
   SIGNAL BU2209_D : STD_LOGIC;
   SIGNAL BU2209_C : STD_LOGIC;
   SIGNAL BU2209_CE : STD_LOGIC;
   SIGNAL BU2209_Q : STD_LOGIC;
   SIGNAL BU2211_D : STD_LOGIC;
   SIGNAL BU2211_C : STD_LOGIC;
   SIGNAL BU2211_CE : STD_LOGIC;
   SIGNAL BU2211_Q : STD_LOGIC;
   SIGNAL BU2213_D : STD_LOGIC;
   SIGNAL BU2213_C : STD_LOGIC;
   SIGNAL BU2213_CE : STD_LOGIC;
   SIGNAL BU2213_Q : STD_LOGIC;
   SIGNAL BU2215_D : STD_LOGIC;
   SIGNAL BU2215_C : STD_LOGIC;
   SIGNAL BU2215_CE : STD_LOGIC;
   SIGNAL BU2215_Q : STD_LOGIC;
   SIGNAL BU2217_D : STD_LOGIC;
   SIGNAL BU2217_C : STD_LOGIC;
   SIGNAL BU2217_CE : STD_LOGIC;
   SIGNAL BU2217_Q : STD_LOGIC;
   SIGNAL BU2219_D : STD_LOGIC;
   SIGNAL BU2219_C : STD_LOGIC;
   SIGNAL BU2219_CE : STD_LOGIC;
   SIGNAL BU2219_Q : STD_LOGIC;
   SIGNAL BU2220_MA : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_MB : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_S : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2220_Q : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_CLK : STD_LOGIC;
   SIGNAL BU2448_D : STD_LOGIC;
   SIGNAL BU2448_C : STD_LOGIC;
   SIGNAL BU2448_CE : STD_LOGIC;
   SIGNAL BU2448_Q : STD_LOGIC;
   SIGNAL BU2452_I0 : STD_LOGIC;
   SIGNAL BU2452_I1 : STD_LOGIC;
   SIGNAL BU2452_I2 : STD_LOGIC;
   SIGNAL BU2452_I3 : STD_LOGIC;
   SIGNAL BU2452_O : STD_LOGIC;
   SIGNAL BU2453_D : STD_LOGIC;
   SIGNAL BU2453_C : STD_LOGIC;
   SIGNAL BU2453_CE : STD_LOGIC;
   SIGNAL BU2453_Q : STD_LOGIC;
   SIGNAL BU2692_DIN : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2692_ND : STD_LOGIC;
   SIGNAL BU2692_RFD : STD_LOGIC;
   SIGNAL BU2692_CLK : STD_LOGIC;
   SIGNAL BU2692_DOUT : STD_LOGIC_VECTOR(46 DOWNTO 0);
   SIGNAL BU2692_RDY : STD_LOGIC;
   SIGNAL BU7718_DIN : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU7718_ND : STD_LOGIC;
   SIGNAL BU7718_RFD : STD_LOGIC;
   SIGNAL BU7718_CLK : STD_LOGIC;
   SIGNAL BU7718_DOUT : STD_LOGIC_VECTOR(46 DOWNTO 0);
   SIGNAL BU7718_RDY : STD_LOGIC;
   SIGNAL BU12513_I0 : STD_LOGIC;
   SIGNAL BU12513_I1 : STD_LOGIC;
   SIGNAL BU12513_I2 : STD_LOGIC;
   SIGNAL BU12513_I3 : STD_LOGIC;
   SIGNAL BU12513_O : STD_LOGIC;
   SIGNAL BU12518_I0 : STD_LOGIC;
   SIGNAL BU12518_I1 : STD_LOGIC;
   SIGNAL BU12518_I2 : STD_LOGIC;
   SIGNAL BU12518_I3 : STD_LOGIC;
   SIGNAL BU12518_O : STD_LOGIC;
   SIGNAL BU12524_D : STD_LOGIC;
   SIGNAL BU12524_CE : STD_LOGIC;
   SIGNAL BU12524_CLK : STD_LOGIC;
   SIGNAL BU12524_A0 : STD_LOGIC;
   SIGNAL BU12524_A1 : STD_LOGIC;
   SIGNAL BU12524_A2 : STD_LOGIC;
   SIGNAL BU12524_A3 : STD_LOGIC;
   SIGNAL BU12524_Q : STD_LOGIC;
   SIGNAL BU12525_D : STD_LOGIC;
   SIGNAL BU12525_CE : STD_LOGIC;
   SIGNAL BU12525_CLK : STD_LOGIC;
   SIGNAL BU12525_A0 : STD_LOGIC;
   SIGNAL BU12525_A1 : STD_LOGIC;
   SIGNAL BU12525_A2 : STD_LOGIC;
   SIGNAL BU12525_A3 : STD_LOGIC;
   SIGNAL BU12525_Q : STD_LOGIC;
   SIGNAL BU12526_D : STD_LOGIC;
   SIGNAL BU12526_CE : STD_LOGIC;
   SIGNAL BU12526_CLK : STD_LOGIC;
   SIGNAL BU12526_A0 : STD_LOGIC;
   SIGNAL BU12526_A1 : STD_LOGIC;
   SIGNAL BU12526_A2 : STD_LOGIC;
   SIGNAL BU12526_A3 : STD_LOGIC;
   SIGNAL BU12526_Q : STD_LOGIC;
   SIGNAL BU12527_D : STD_LOGIC;
   SIGNAL BU12527_CE : STD_LOGIC;
   SIGNAL BU12527_CLK : STD_LOGIC;
   SIGNAL BU12527_A0 : STD_LOGIC;
   SIGNAL BU12527_A1 : STD_LOGIC;
   SIGNAL BU12527_A2 : STD_LOGIC;
   SIGNAL BU12527_A3 : STD_LOGIC;
   SIGNAL BU12527_Q : STD_LOGIC;
   SIGNAL BU12528_D : STD_LOGIC;
   SIGNAL BU12528_CE : STD_LOGIC;
   SIGNAL BU12528_CLK : STD_LOGIC;
   SIGNAL BU12528_A0 : STD_LOGIC;
   SIGNAL BU12528_A1 : STD_LOGIC;
   SIGNAL BU12528_A2 : STD_LOGIC;
   SIGNAL BU12528_A3 : STD_LOGIC;
   SIGNAL BU12528_Q : STD_LOGIC;
   SIGNAL BU12529_D : STD_LOGIC;
   SIGNAL BU12529_CE : STD_LOGIC;
   SIGNAL BU12529_CLK : STD_LOGIC;
   SIGNAL BU12529_A0 : STD_LOGIC;
   SIGNAL BU12529_A1 : STD_LOGIC;
   SIGNAL BU12529_A2 : STD_LOGIC;
   SIGNAL BU12529_A3 : STD_LOGIC;
   SIGNAL BU12529_Q : STD_LOGIC;
   SIGNAL BU12530_D : STD_LOGIC;
   SIGNAL BU12530_CE : STD_LOGIC;
   SIGNAL BU12530_CLK : STD_LOGIC;
   SIGNAL BU12530_A0 : STD_LOGIC;
   SIGNAL BU12530_A1 : STD_LOGIC;
   SIGNAL BU12530_A2 : STD_LOGIC;
   SIGNAL BU12530_A3 : STD_LOGIC;
   SIGNAL BU12530_Q : STD_LOGIC;
   SIGNAL BU12531_D : STD_LOGIC;
   SIGNAL BU12531_CE : STD_LOGIC;
   SIGNAL BU12531_CLK : STD_LOGIC;
   SIGNAL BU12531_A0 : STD_LOGIC;
   SIGNAL BU12531_A1 : STD_LOGIC;
   SIGNAL BU12531_A2 : STD_LOGIC;
   SIGNAL BU12531_A3 : STD_LOGIC;
   SIGNAL BU12531_Q : STD_LOGIC;
   SIGNAL BU12532_D : STD_LOGIC;
   SIGNAL BU12532_CE : STD_LOGIC;
   SIGNAL BU12532_CLK : STD_LOGIC;
   SIGNAL BU12532_A0 : STD_LOGIC;
   SIGNAL BU12532_A1 : STD_LOGIC;
   SIGNAL BU12532_A2 : STD_LOGIC;
   SIGNAL BU12532_A3 : STD_LOGIC;
   SIGNAL BU12532_Q : STD_LOGIC;
   SIGNAL BU12533_D : STD_LOGIC;
   SIGNAL BU12533_CE : STD_LOGIC;
   SIGNAL BU12533_CLK : STD_LOGIC;
   SIGNAL BU12533_A0 : STD_LOGIC;
   SIGNAL BU12533_A1 : STD_LOGIC;
   SIGNAL BU12533_A2 : STD_LOGIC;
   SIGNAL BU12533_A3 : STD_LOGIC;
   SIGNAL BU12533_Q : STD_LOGIC;
   SIGNAL BU12534_D : STD_LOGIC;
   SIGNAL BU12534_CE : STD_LOGIC;
   SIGNAL BU12534_CLK : STD_LOGIC;
   SIGNAL BU12534_A0 : STD_LOGIC;
   SIGNAL BU12534_A1 : STD_LOGIC;
   SIGNAL BU12534_A2 : STD_LOGIC;
   SIGNAL BU12534_A3 : STD_LOGIC;
   SIGNAL BU12534_Q : STD_LOGIC;
   SIGNAL BU12535_D : STD_LOGIC;
   SIGNAL BU12535_CE : STD_LOGIC;
   SIGNAL BU12535_CLK : STD_LOGIC;
   SIGNAL BU12535_A0 : STD_LOGIC;
   SIGNAL BU12535_A1 : STD_LOGIC;
   SIGNAL BU12535_A2 : STD_LOGIC;
   SIGNAL BU12535_A3 : STD_LOGIC;
   SIGNAL BU12535_Q : STD_LOGIC;
   SIGNAL BU12536_D : STD_LOGIC;
   SIGNAL BU12536_CE : STD_LOGIC;
   SIGNAL BU12536_CLK : STD_LOGIC;
   SIGNAL BU12536_A0 : STD_LOGIC;
   SIGNAL BU12536_A1 : STD_LOGIC;
   SIGNAL BU12536_A2 : STD_LOGIC;
   SIGNAL BU12536_A3 : STD_LOGIC;
   SIGNAL BU12536_Q : STD_LOGIC;
   SIGNAL BU12537_D : STD_LOGIC;
   SIGNAL BU12537_CE : STD_LOGIC;
   SIGNAL BU12537_CLK : STD_LOGIC;
   SIGNAL BU12537_A0 : STD_LOGIC;
   SIGNAL BU12537_A1 : STD_LOGIC;
   SIGNAL BU12537_A2 : STD_LOGIC;
   SIGNAL BU12537_A3 : STD_LOGIC;
   SIGNAL BU12537_Q : STD_LOGIC;
   SIGNAL BU12538_D : STD_LOGIC;
   SIGNAL BU12538_CE : STD_LOGIC;
   SIGNAL BU12538_CLK : STD_LOGIC;
   SIGNAL BU12538_A0 : STD_LOGIC;
   SIGNAL BU12538_A1 : STD_LOGIC;
   SIGNAL BU12538_A2 : STD_LOGIC;
   SIGNAL BU12538_A3 : STD_LOGIC;
   SIGNAL BU12538_Q : STD_LOGIC;
   SIGNAL BU12539_D : STD_LOGIC;
   SIGNAL BU12539_CE : STD_LOGIC;
   SIGNAL BU12539_CLK : STD_LOGIC;
   SIGNAL BU12539_A0 : STD_LOGIC;
   SIGNAL BU12539_A1 : STD_LOGIC;
   SIGNAL BU12539_A2 : STD_LOGIC;
   SIGNAL BU12539_A3 : STD_LOGIC;
   SIGNAL BU12539_Q : STD_LOGIC;
   SIGNAL BU12540_D : STD_LOGIC;
   SIGNAL BU12540_CE : STD_LOGIC;
   SIGNAL BU12540_CLK : STD_LOGIC;
   SIGNAL BU12540_A0 : STD_LOGIC;
   SIGNAL BU12540_A1 : STD_LOGIC;
   SIGNAL BU12540_A2 : STD_LOGIC;
   SIGNAL BU12540_A3 : STD_LOGIC;
   SIGNAL BU12540_Q : STD_LOGIC;
   SIGNAL BU12541_D : STD_LOGIC;
   SIGNAL BU12541_CE : STD_LOGIC;
   SIGNAL BU12541_CLK : STD_LOGIC;
   SIGNAL BU12541_A0 : STD_LOGIC;
   SIGNAL BU12541_A1 : STD_LOGIC;
   SIGNAL BU12541_A2 : STD_LOGIC;
   SIGNAL BU12541_A3 : STD_LOGIC;
   SIGNAL BU12541_Q : STD_LOGIC;
   SIGNAL BU12542_D : STD_LOGIC;
   SIGNAL BU12542_CE : STD_LOGIC;
   SIGNAL BU12542_CLK : STD_LOGIC;
   SIGNAL BU12542_A0 : STD_LOGIC;
   SIGNAL BU12542_A1 : STD_LOGIC;
   SIGNAL BU12542_A2 : STD_LOGIC;
   SIGNAL BU12542_A3 : STD_LOGIC;
   SIGNAL BU12542_Q : STD_LOGIC;
   SIGNAL BU12543_D : STD_LOGIC;
   SIGNAL BU12543_CE : STD_LOGIC;
   SIGNAL BU12543_CLK : STD_LOGIC;
   SIGNAL BU12543_A0 : STD_LOGIC;
   SIGNAL BU12543_A1 : STD_LOGIC;
   SIGNAL BU12543_A2 : STD_LOGIC;
   SIGNAL BU12543_A3 : STD_LOGIC;
   SIGNAL BU12543_Q : STD_LOGIC;
   SIGNAL BU12544_D : STD_LOGIC;
   SIGNAL BU12544_CE : STD_LOGIC;
   SIGNAL BU12544_CLK : STD_LOGIC;
   SIGNAL BU12544_A0 : STD_LOGIC;
   SIGNAL BU12544_A1 : STD_LOGIC;
   SIGNAL BU12544_A2 : STD_LOGIC;
   SIGNAL BU12544_A3 : STD_LOGIC;
   SIGNAL BU12544_Q : STD_LOGIC;
   SIGNAL BU12545_D : STD_LOGIC;
   SIGNAL BU12545_CE : STD_LOGIC;
   SIGNAL BU12545_CLK : STD_LOGIC;
   SIGNAL BU12545_A0 : STD_LOGIC;
   SIGNAL BU12545_A1 : STD_LOGIC;
   SIGNAL BU12545_A2 : STD_LOGIC;
   SIGNAL BU12545_A3 : STD_LOGIC;
   SIGNAL BU12545_Q : STD_LOGIC;
   SIGNAL BU12546_D : STD_LOGIC;
   SIGNAL BU12546_CE : STD_LOGIC;
   SIGNAL BU12546_CLK : STD_LOGIC;
   SIGNAL BU12546_A0 : STD_LOGIC;
   SIGNAL BU12546_A1 : STD_LOGIC;
   SIGNAL BU12546_A2 : STD_LOGIC;
   SIGNAL BU12546_A3 : STD_LOGIC;
   SIGNAL BU12546_Q : STD_LOGIC;
   SIGNAL BU12547_D : STD_LOGIC;
   SIGNAL BU12547_CE : STD_LOGIC;
   SIGNAL BU12547_CLK : STD_LOGIC;
   SIGNAL BU12547_A0 : STD_LOGIC;
   SIGNAL BU12547_A1 : STD_LOGIC;
   SIGNAL BU12547_A2 : STD_LOGIC;
   SIGNAL BU12547_A3 : STD_LOGIC;
   SIGNAL BU12547_Q : STD_LOGIC;
   SIGNAL BU12548_D : STD_LOGIC;
   SIGNAL BU12548_CE : STD_LOGIC;
   SIGNAL BU12548_CLK : STD_LOGIC;
   SIGNAL BU12548_A0 : STD_LOGIC;
   SIGNAL BU12548_A1 : STD_LOGIC;
   SIGNAL BU12548_A2 : STD_LOGIC;
   SIGNAL BU12548_A3 : STD_LOGIC;
   SIGNAL BU12548_Q : STD_LOGIC;
   SIGNAL BU12549_D : STD_LOGIC;
   SIGNAL BU12549_CE : STD_LOGIC;
   SIGNAL BU12549_CLK : STD_LOGIC;
   SIGNAL BU12549_A0 : STD_LOGIC;
   SIGNAL BU12549_A1 : STD_LOGIC;
   SIGNAL BU12549_A2 : STD_LOGIC;
   SIGNAL BU12549_A3 : STD_LOGIC;
   SIGNAL BU12549_Q : STD_LOGIC;
   SIGNAL BU12550_Q : STD_LOGIC_VECTOR(3 DOWNTO 0);
   SIGNAL BU12550_CLK : STD_LOGIC;
   SIGNAL BU12550_UP : STD_LOGIC;
   SIGNAL BU12550_CE : STD_LOGIC;
   SIGNAL BU12579_I0 : STD_LOGIC;
   SIGNAL BU12579_I1 : STD_LOGIC;
   SIGNAL BU12579_I2 : STD_LOGIC;
   SIGNAL BU12579_I3 : STD_LOGIC;
   SIGNAL BU12579_O : STD_LOGIC;
   SIGNAL BU12583_I0 : STD_LOGIC;
   SIGNAL BU12583_I1 : STD_LOGIC;
   SIGNAL BU12583_I2 : STD_LOGIC;
   SIGNAL BU12583_I3 : STD_LOGIC;
   SIGNAL BU12583_O : STD_LOGIC;
   SIGNAL BU12584_D : STD_LOGIC;
   SIGNAL BU12584_C : STD_LOGIC;
   SIGNAL BU12584_CE : STD_LOGIC;
   SIGNAL BU12584_Q : STD_LOGIC;
   SIGNAL BU12587_I0 : STD_LOGIC;
   SIGNAL BU12587_I1 : STD_LOGIC;
   SIGNAL BU12587_I2 : STD_LOGIC;
   SIGNAL BU12587_I3 : STD_LOGIC;
   SIGNAL BU12587_O : STD_LOGIC;
   SIGNAL BU12588_ND : STD_LOGIC;
   SIGNAL BU12588_RDY : STD_LOGIC;
   SIGNAL BU12588_CLK : STD_LOGIC;
   SIGNAL BU12588_RFD : STD_LOGIC;
   SIGNAL BU12588_DIN : STD_LOGIC_VECTOR(25 DOWNTO 0);
   SIGNAL BU12588_DOUT : STD_LOGIC_VECTOR(42 DOWNTO 0);
   SIGNAL BU19118_I : STD_LOGIC_VECTOR(26 DOWNTO 0);
   SIGNAL BU19118_O : STD_LOGIC;
   SIGNAL BU19149_I0 : STD_LOGIC;
   SIGNAL BU19149_I1 : STD_LOGIC;
   SIGNAL BU19149_I2 : STD_LOGIC;
   SIGNAL BU19149_I3 : STD_LOGIC;
   SIGNAL BU19149_O : STD_LOGIC;
   SIGNAL BU19150_A : STD_LOGIC_VECTOR(15 DOWNTO 0);
   SIGNAL BU19150_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU19150_S : STD_LOGIC_VECTOR(16 DOWNTO 0);
   SIGNAL BU19219_I0 : STD_LOGIC;
   SIGNAL BU19219_I1 : STD_LOGIC;
   SIGNAL BU19219_I2 : STD_LOGIC;
   SIGNAL BU19219_I3 : STD_LOGIC;
   SIGNAL BU19219_O : STD_LOGIC;
   SIGNAL BU19221_I0 : STD_LOGIC;
   SIGNAL BU19221_I1 : STD_LOGIC;
   SIGNAL BU19221_I2 : STD_LOGIC;
   SIGNAL BU19221_I3 : STD_LOGIC;
   SIGNAL BU19221_O : STD_LOGIC;
   SIGNAL BU19222_D : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU19222_Q : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU19222_CLK : STD_LOGIC;
   SIGNAL BU19222_SCLR : STD_LOGIC;
   SIGNAL BU19222_SSET : STD_LOGIC;
   SIGNAL BU19283_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU19283_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU19283_CLK : STD_LOGIC;
   SIGNAL BU19283_SCLR : STD_LOGIC;
   SIGNAL BU19283_SSET : STD_LOGIC;
   SIGNAL BU19290_D : STD_LOGIC;
   SIGNAL BU19290_C : STD_LOGIC;
   SIGNAL BU19290_CE : STD_LOGIC;
   SIGNAL BU19290_Q : STD_LOGIC;
   SIGNAL BU19293_ND : STD_LOGIC;
   SIGNAL BU19293_RDY : STD_LOGIC;
   SIGNAL BU19293_CLK : STD_LOGIC;
   SIGNAL BU19293_RFD : STD_LOGIC;
   SIGNAL BU19293_DIN : STD_LOGIC_VECTOR(15 DOWNTO 0);
   SIGNAL BU19293_SEL_O : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU19293_DOUT : STD_LOGIC_VECTOR(34 DOWNTO 0);
   SIGNAL BU22774_I0 : STD_LOGIC;
   SIGNAL BU22774_I1 : STD_LOGIC;
   SIGNAL BU22774_I2 : STD_LOGIC;
   SIGNAL BU22774_I3 : STD_LOGIC;
   SIGNAL BU22774_O : STD_LOGIC;
   SIGNAL BU22776_I0 : STD_LOGIC;
   SIGNAL BU22776_I1 : STD_LOGIC;
   SIGNAL BU22776_I2 : STD_LOGIC;
   SIGNAL BU22776_I3 : STD_LOGIC;
   SIGNAL BU22776_O : STD_LOGIC;
   SIGNAL BU22779_D : STD_LOGIC;
   SIGNAL BU22779_C : STD_LOGIC;
   SIGNAL BU22779_CE : STD_LOGIC;
   SIGNAL BU22779_Q : STD_LOGIC;
   SIGNAL BU22784_I : STD_LOGIC_VECTOR(4 DOWNTO 0);
   SIGNAL BU22784_O : STD_LOGIC;
   SIGNAL BU22793_I0 : STD_LOGIC;
   SIGNAL BU22793_I1 : STD_LOGIC;
   SIGNAL BU22793_I2 : STD_LOGIC;
   SIGNAL BU22793_I3 : STD_LOGIC;
   SIGNAL BU22793_O : STD_LOGIC;
   SIGNAL BU22794_A : STD_LOGIC_VECTOR(29 DOWNTO 0);
   SIGNAL BU22794_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU22794_S : STD_LOGIC_VECTOR(30 DOWNTO 0);
   SIGNAL BU22919_I0 : STD_LOGIC;
   SIGNAL BU22919_I1 : STD_LOGIC;
   SIGNAL BU22919_I2 : STD_LOGIC;
   SIGNAL BU22919_I3 : STD_LOGIC;
   SIGNAL BU22919_O : STD_LOGIC;
   SIGNAL BU22921_I0 : STD_LOGIC;
   SIGNAL BU22921_I1 : STD_LOGIC;
   SIGNAL BU22921_I2 : STD_LOGIC;
   SIGNAL BU22921_I3 : STD_LOGIC;
   SIGNAL BU22921_O : STD_LOGIC;
   SIGNAL BU22922_D : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU22922_Q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU22922_CLK : STD_LOGIC;
   SIGNAL BU22922_CE : STD_LOGIC;
   SIGNAL BU22922_SCLR : STD_LOGIC;
   SIGNAL BU22922_SSET : STD_LOGIC;
   SIGNAL BU23042_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU23042_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU23042_CLK : STD_LOGIC;
   SIGNAL BU23042_CE : STD_LOGIC;
   SIGNAL BU23042_SCLR : STD_LOGIC;
   SIGNAL BU23042_SSET : STD_LOGIC;
   SIGNAL BU23054_I : STD_LOGIC_VECTOR(4 DOWNTO 0);
   SIGNAL BU23054_O : STD_LOGIC;
   SIGNAL BU23063_I0 : STD_LOGIC;
   SIGNAL BU23063_I1 : STD_LOGIC;
   SIGNAL BU23063_I2 : STD_LOGIC;
   SIGNAL BU23063_I3 : STD_LOGIC;
   SIGNAL BU23063_O : STD_LOGIC;
   SIGNAL BU23064_A : STD_LOGIC_VECTOR(29 DOWNTO 0);
   SIGNAL BU23064_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU23064_S : STD_LOGIC_VECTOR(30 DOWNTO 0);
   SIGNAL BU23189_I0 : STD_LOGIC;
   SIGNAL BU23189_I1 : STD_LOGIC;
   SIGNAL BU23189_I2 : STD_LOGIC;
   SIGNAL BU23189_I3 : STD_LOGIC;
   SIGNAL BU23189_O : STD_LOGIC;
   SIGNAL BU23191_I0 : STD_LOGIC;
   SIGNAL BU23191_I1 : STD_LOGIC;
   SIGNAL BU23191_I2 : STD_LOGIC;
   SIGNAL BU23191_I3 : STD_LOGIC;
   SIGNAL BU23191_O : STD_LOGIC;
   SIGNAL BU23192_D : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU23192_Q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU23192_CLK : STD_LOGIC;
   SIGNAL BU23192_CE : STD_LOGIC;
   SIGNAL BU23192_SCLR : STD_LOGIC;
   SIGNAL BU23192_SSET : STD_LOGIC;
   SIGNAL BU23312_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU23312_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU23312_CLK : STD_LOGIC;
   SIGNAL BU23312_CE : STD_LOGIC;
   SIGNAL BU23312_SCLR : STD_LOGIC;
   SIGNAL BU23312_SSET : STD_LOGIC;
   SIGNAL n0 : STD_LOGIC := '0';
   SIGNAL n1 : STD_LOGIC := '1';
   SIGNAL n2 : STD_LOGIC;
   SIGNAL n3 : STD_LOGIC;
   SIGNAL n4 : STD_LOGIC;
   SIGNAL n5 : STD_LOGIC;
   SIGNAL n6 : STD_LOGIC;
   SIGNAL n7 : STD_LOGIC;
   SIGNAL n8 : STD_LOGIC;
   SIGNAL n9 : STD_LOGIC;
   SIGNAL n10 : STD_LOGIC;
   SIGNAL n11 : STD_LOGIC;
   SIGNAL n12 : STD_LOGIC;
   SIGNAL n13 : STD_LOGIC;
   SIGNAL n14 : STD_LOGIC;
   SIGNAL n15 : STD_LOGIC;
   SIGNAL n16 : STD_LOGIC;
   SIGNAL n17 : STD_LOGIC;
   SIGNAL n18 : STD_LOGIC;
   SIGNAL n19 : STD_LOGIC;
   SIGNAL n20 : STD_LOGIC;
   SIGNAL n21 : STD_LOGIC;
   SIGNAL n22 : STD_LOGIC;
   SIGNAL n23 : STD_LOGIC;
   SIGNAL n24 : STD_LOGIC;
   SIGNAL n25 : STD_LOGIC;
   SIGNAL n26 : STD_LOGIC;
   SIGNAL n27 : STD_LOGIC;
   SIGNAL n28 : STD_LOGIC;
   SIGNAL n29 : STD_LOGIC;
   SIGNAL n30 : STD_LOGIC;
   SIGNAL n31 : STD_LOGIC;
   SIGNAL n32 : STD_LOGIC;
   SIGNAL n33 : STD_LOGIC;
   SIGNAL n34 : STD_LOGIC;
   SIGNAL n35 : STD_LOGIC;
   SIGNAL n36 : STD_LOGIC;
   SIGNAL n37 : STD_LOGIC;
   SIGNAL n38 : STD_LOGIC;
   SIGNAL n39 : STD_LOGIC;
   SIGNAL n40 : STD_LOGIC;
   SIGNAL n41 : STD_LOGIC;
   SIGNAL n42 : STD_LOGIC;
   SIGNAL n43 : STD_LOGIC;
   SIGNAL n44 : STD_LOGIC;
   SIGNAL n45 : STD_LOGIC;
   SIGNAL n46 : STD_LOGIC;
   SIGNAL n47 : STD_LOGIC;
   SIGNAL n48 : STD_LOGIC;
   SIGNAL n49 : STD_LOGIC;
   SIGNAL n50 : STD_LOGIC;
   SIGNAL n54 : STD_LOGIC;
   SIGNAL n55 : STD_LOGIC;
   SIGNAL n58 : STD_LOGIC;
   SIGNAL n59 : STD_LOGIC;
   SIGNAL n60 : STD_LOGIC;
   SIGNAL n61 : STD_LOGIC;
   SIGNAL n62 : STD_LOGIC;
   SIGNAL n63 : STD_LOGIC;
   SIGNAL n64 : STD_LOGIC;
   SIGNAL n65 : STD_LOGIC;
   SIGNAL n66 : STD_LOGIC;
   SIGNAL n67 : STD_LOGIC;
   SIGNAL n68 : STD_LOGIC;
   SIGNAL n69 : STD_LOGIC;
   SIGNAL n70 : STD_LOGIC;
   SIGNAL n71 : STD_LOGIC;
   SIGNAL n72 : STD_LOGIC;
   SIGNAL n73 : STD_LOGIC;
   SIGNAL n74 : STD_LOGIC;
   SIGNAL n75 : STD_LOGIC;
   SIGNAL n76 : STD_LOGIC;
   SIGNAL n77 : STD_LOGIC;
   SIGNAL n78 : STD_LOGIC;
   SIGNAL n79 : STD_LOGIC;
   SIGNAL n80 : STD_LOGIC;
   SIGNAL n81 : STD_LOGIC;
   SIGNAL n82 : STD_LOGIC;
   SIGNAL n83 : STD_LOGIC;
   SIGNAL n84 : STD_LOGIC;
   SIGNAL n85 : STD_LOGIC;
   SIGNAL n86 : STD_LOGIC;
   SIGNAL n87 : STD_LOGIC;
   SIGNAL n88 : STD_LOGIC;
   SIGNAL n89 : STD_LOGIC;
   SIGNAL n90 : STD_LOGIC;
   SIGNAL n91 : STD_LOGIC;
   SIGNAL n92 : STD_LOGIC;
   SIGNAL n93 : STD_LOGIC;
   SIGNAL n94 : STD_LOGIC;
   SIGNAL n95 : STD_LOGIC;
   SIGNAL n96 : STD_LOGIC;
   SIGNAL n97 : STD_LOGIC;
   SIGNAL n98 : STD_LOGIC;
   SIGNAL n99 : STD_LOGIC;
   SIGNAL n100 : STD_LOGIC;
   SIGNAL n101 : STD_LOGIC;
   SIGNAL n102 : STD_LOGIC;
   SIGNAL n103 : STD_LOGIC;
   SIGNAL n104 : STD_LOGIC;
   SIGNAL n105 : STD_LOGIC;
   SIGNAL n106 : STD_LOGIC;
   SIGNAL n107 : STD_LOGIC;
   SIGNAL n108 : STD_LOGIC;
   SIGNAL n109 : STD_LOGIC;
   SIGNAL n110 : STD_LOGIC;
   SIGNAL n111 : STD_LOGIC;
   SIGNAL n112 : STD_LOGIC;
   SIGNAL n113 : STD_LOGIC;
   SIGNAL n114 : STD_LOGIC;
   SIGNAL n115 : STD_LOGIC;
   SIGNAL n116 : STD_LOGIC;
   SIGNAL n117 : STD_LOGIC;
   SIGNAL n118 : STD_LOGIC;
   SIGNAL n119 : STD_LOGIC;
   SIGNAL n120 : STD_LOGIC;
   SIGNAL n121 : STD_LOGIC;
   SIGNAL n122 : STD_LOGIC;
   SIGNAL n123 : STD_LOGIC;
   SIGNAL n124 : STD_LOGIC;
   SIGNAL n125 : STD_LOGIC;
   SIGNAL n126 : STD_LOGIC;
   SIGNAL n127 : STD_LOGIC;
   SIGNAL n128 : STD_LOGIC;
   SIGNAL n129 : STD_LOGIC;
   SIGNAL n130 : STD_LOGIC;
   SIGNAL n131 : STD_LOGIC;
   SIGNAL n132 : STD_LOGIC;
   SIGNAL n133 : STD_LOGIC;
   SIGNAL n134 : STD_LOGIC;
   SIGNAL n135 : STD_LOGIC;
   SIGNAL n136 : STD_LOGIC;
   SIGNAL n137 : STD_LOGIC;
   SIGNAL n138 : STD_LOGIC;
   SIGNAL n139 : STD_LOGIC;
   SIGNAL n140 : STD_LOGIC;
   SIGNAL n141 : STD_LOGIC;
   SIGNAL n142 : STD_LOGIC;
   SIGNAL n143 : STD_LOGIC;
   SIGNAL n144 : STD_LOGIC;
   SIGNAL n145 : STD_LOGIC;
   SIGNAL n146 : STD_LOGIC;
   SIGNAL n147 : STD_LOGIC;
   SIGNAL n148 : STD_LOGIC;
   SIGNAL n149 : STD_LOGIC;
   SIGNAL n150 : STD_LOGIC;
   SIGNAL n151 : STD_LOGIC;
   SIGNAL n152 : STD_LOGIC;
   SIGNAL n153 : STD_LOGIC;
   SIGNAL n154 : STD_LOGIC;
   SIGNAL n155 : STD_LOGIC;
   SIGNAL n156 : STD_LOGIC;
   SIGNAL n157 : STD_LOGIC;
   SIGNAL n158 : STD_LOGIC;
   SIGNAL n159 : STD_LOGIC;
   SIGNAL n160 : STD_LOGIC;
   SIGNAL n161 : STD_LOGIC;
   SIGNAL n162 : STD_LOGIC;
   SIGNAL n163 : STD_LOGIC;
   SIGNAL n164 : STD_LOGIC;
   SIGNAL n165 : STD_LOGIC;
   SIGNAL n166 : STD_LOGIC;
   SIGNAL n167 : STD_LOGIC;
   SIGNAL n168 : STD_LOGIC;
   SIGNAL n169 : STD_LOGIC;
   SIGNAL n170 : STD_LOGIC;
   SIGNAL n171 : STD_LOGIC;
   SIGNAL n172 : STD_LOGIC;
   SIGNAL n173 : STD_LOGIC;
   SIGNAL n174 : STD_LOGIC;
   SIGNAL n175 : STD_LOGIC;
   SIGNAL n176 : STD_LOGIC;
   SIGNAL n177 : STD_LOGIC;
   SIGNAL n178 : STD_LOGIC;
   SIGNAL n179 : STD_LOGIC;
   SIGNAL n180 : STD_LOGIC;
   SIGNAL n181 : STD_LOGIC;
   SIGNAL n182 : STD_LOGIC;
   SIGNAL n183 : STD_LOGIC;
   SIGNAL n184 : STD_LOGIC;
   SIGNAL n185 : STD_LOGIC;
   SIGNAL n186 : STD_LOGIC;
   SIGNAL n187 : STD_LOGIC;
   SIGNAL n188 : STD_LOGIC;
   SIGNAL n189 : STD_LOGIC;
   SIGNAL n190 : STD_LOGIC;
   SIGNAL n191 : STD_LOGIC;
   SIGNAL n192 : STD_LOGIC;
   SIGNAL n193 : STD_LOGIC;
   SIGNAL n194 : STD_LOGIC;
   SIGNAL n195 : STD_LOGIC;
   SIGNAL n196 : STD_LOGIC;
   SIGNAL n197 : STD_LOGIC;
   SIGNAL n198 : STD_LOGIC;
   SIGNAL n199 : STD_LOGIC;
   SIGNAL n200 : STD_LOGIC;
   SIGNAL n201 : STD_LOGIC;
   SIGNAL n202 : STD_LOGIC;
   SIGNAL n203 : STD_LOGIC;
   SIGNAL n204 : STD_LOGIC;
   SIGNAL n205 : STD_LOGIC;
   SIGNAL n206 : STD_LOGIC;
   SIGNAL n207 : STD_LOGIC;
   SIGNAL n208 : STD_LOGIC;
   SIGNAL n209 : STD_LOGIC;
   SIGNAL n210 : STD_LOGIC;
   SIGNAL n211 : STD_LOGIC;
   SIGNAL n212 : STD_LOGIC;
   SIGNAL n213 : STD_LOGIC;
   SIGNAL n214 : STD_LOGIC;
   SIGNAL n215 : STD_LOGIC;
   SIGNAL n216 : STD_LOGIC;
   SIGNAL n217 : STD_LOGIC;
   SIGNAL n218 : STD_LOGIC;
   SIGNAL n219 : STD_LOGIC;
   SIGNAL n220 : STD_LOGIC;
   SIGNAL n221 : STD_LOGIC;
   SIGNAL n222 : STD_LOGIC;
   SIGNAL n223 : STD_LOGIC;
   SIGNAL n224 : STD_LOGIC;
   SIGNAL n225 : STD_LOGIC;
   SIGNAL n226 : STD_LOGIC;
   SIGNAL n227 : STD_LOGIC;
   SIGNAL n228 : STD_LOGIC;
   SIGNAL n229 : STD_LOGIC;
   SIGNAL n230 : STD_LOGIC;
   SIGNAL n231 : STD_LOGIC;
   SIGNAL n232 : STD_LOGIC;
   SIGNAL n233 : STD_LOGIC;
   SIGNAL n234 : STD_LOGIC;
   SIGNAL n235 : STD_LOGIC;
   SIGNAL n236 : STD_LOGIC;
   SIGNAL n237 : STD_LOGIC;
   SIGNAL n238 : STD_LOGIC;
   SIGNAL n239 : STD_LOGIC;
   SIGNAL n240 : STD_LOGIC;
   SIGNAL n241 : STD_LOGIC;
   SIGNAL n242 : STD_LOGIC;
   SIGNAL n243 : STD_LOGIC;
   SIGNAL n244 : STD_LOGIC;
   SIGNAL n245 : STD_LOGIC;
   SIGNAL n246 : STD_LOGIC;
   SIGNAL n247 : STD_LOGIC;
   SIGNAL n248 : STD_LOGIC;
   SIGNAL n249 : STD_LOGIC;
   SIGNAL n250 : STD_LOGIC;
   SIGNAL n251 : STD_LOGIC;
   SIGNAL n252 : STD_LOGIC;
   SIGNAL n253 : STD_LOGIC;
   SIGNAL n254 : STD_LOGIC;
   SIGNAL n294 : STD_LOGIC;
   SIGNAL n341 : STD_LOGIC;
   SIGNAL n342 : STD_LOGIC;
   SIGNAL n343 : STD_LOGIC;
   SIGNAL n415 : STD_LOGIC;
   SIGNAL n416 : STD_LOGIC;
   SIGNAL n417 : STD_LOGIC;
   SIGNAL n418 : STD_LOGIC;
   SIGNAL n419 : STD_LOGIC;
   SIGNAL n420 : STD_LOGIC;
   SIGNAL n421 : STD_LOGIC;
   SIGNAL n422 : STD_LOGIC;
   SIGNAL n423 : STD_LOGIC;
   SIGNAL n424 : STD_LOGIC;
   SIGNAL n425 : STD_LOGIC;
   SIGNAL n426 : STD_LOGIC;
   SIGNAL n427 : STD_LOGIC;
   SIGNAL n428 : STD_LOGIC;
   SIGNAL n429 : STD_LOGIC;
   SIGNAL n460 : STD_LOGIC;
   SIGNAL n461 : STD_LOGIC;
   SIGNAL n462 : STD_LOGIC;
   SIGNAL n463 : STD_LOGIC;
   SIGNAL n464 : STD_LOGIC;
   SIGNAL n465 : STD_LOGIC;
   SIGNAL n466 : STD_LOGIC;
   SIGNAL n467 : STD_LOGIC;
   SIGNAL n468 : STD_LOGIC;
   SIGNAL n469 : STD_LOGIC;
   SIGNAL n470 : STD_LOGIC;
   SIGNAL n471 : STD_LOGIC;
   SIGNAL n472 : STD_LOGIC;
   SIGNAL n473 : STD_LOGIC;
   SIGNAL n474 : STD_LOGIC;
   SIGNAL n475 : STD_LOGIC;
   SIGNAL n476 : STD_LOGIC;
   SIGNAL n477 : STD_LOGIC;
   SIGNAL n478 : STD_LOGIC;
   SIGNAL n479 : STD_LOGIC;
   SIGNAL n480 : STD_LOGIC;
   SIGNAL n481 : STD_LOGIC;
   SIGNAL n482 : STD_LOGIC;
   SIGNAL n483 : STD_LOGIC;
   SIGNAL n484 : STD_LOGIC;
   SIGNAL n485 : STD_LOGIC;
   SIGNAL n486 : STD_LOGIC;
   SIGNAL n487 : STD_LOGIC;
   SIGNAL n488 : STD_LOGIC;
   SIGNAL n547 : STD_LOGIC;
   SIGNAL n577 : STD_LOGIC;
   SIGNAL n578 : STD_LOGIC;
   SIGNAL n579 : STD_LOGIC;
   SIGNAL n580 : STD_LOGIC;
   SIGNAL n581 : STD_LOGIC;
   SIGNAL n582 : STD_LOGIC;
   SIGNAL n583 : STD_LOGIC;
   SIGNAL n584 : STD_LOGIC;
   SIGNAL n585 : STD_LOGIC;
   SIGNAL n586 : STD_LOGIC;
   SIGNAL n587 : STD_LOGIC;
   SIGNAL n588 : STD_LOGIC;
   SIGNAL n589 : STD_LOGIC;
   SIGNAL n590 : STD_LOGIC;
   SIGNAL n619 : STD_LOGIC;
   SIGNAL n620 : STD_LOGIC;
   SIGNAL n621 : STD_LOGIC;
   SIGNAL n622 : STD_LOGIC;
   SIGNAL n623 : STD_LOGIC;
   SIGNAL n624 : STD_LOGIC;
   SIGNAL n625 : STD_LOGIC;
   SIGNAL n626 : STD_LOGIC;
   SIGNAL n627 : STD_LOGIC;
   SIGNAL n628 : STD_LOGIC;
   SIGNAL n629 : STD_LOGIC;
   SIGNAL n630 : STD_LOGIC;
   SIGNAL n631 : STD_LOGIC;
   SIGNAL n632 : STD_LOGIC;
   SIGNAL n633 : STD_LOGIC;
   SIGNAL n664 : STD_LOGIC;
   SIGNAL n665 : STD_LOGIC;
   SIGNAL n666 : STD_LOGIC;
   SIGNAL n667 : STD_LOGIC;
   SIGNAL n668 : STD_LOGIC;
   SIGNAL n669 : STD_LOGIC;
   SIGNAL n670 : STD_LOGIC;
   SIGNAL n671 : STD_LOGIC;
   SIGNAL n672 : STD_LOGIC;
   SIGNAL n673 : STD_LOGIC;
   SIGNAL n674 : STD_LOGIC;
   SIGNAL n675 : STD_LOGIC;
   SIGNAL n676 : STD_LOGIC;
   SIGNAL n677 : STD_LOGIC;
   SIGNAL n678 : STD_LOGIC;
   SIGNAL n679 : STD_LOGIC;
   SIGNAL n680 : STD_LOGIC;
   SIGNAL n681 : STD_LOGIC;
   SIGNAL n682 : STD_LOGIC;
   SIGNAL n683 : STD_LOGIC;
   SIGNAL n684 : STD_LOGIC;
   SIGNAL n685 : STD_LOGIC;
   SIGNAL n686 : STD_LOGIC;
   SIGNAL n687 : STD_LOGIC;
   SIGNAL n688 : STD_LOGIC;
   SIGNAL n689 : STD_LOGIC;
   SIGNAL n690 : STD_LOGIC;
   SIGNAL n691 : STD_LOGIC;
   SIGNAL n692 : STD_LOGIC;
   SIGNAL n927 : STD_LOGIC;
   SIGNAL n928 : STD_LOGIC;
   SIGNAL n929 : STD_LOGIC;
   SIGNAL n930 : STD_LOGIC;
   SIGNAL n931 : STD_LOGIC;
   SIGNAL n932 : STD_LOGIC;
   SIGNAL n933 : STD_LOGIC;
   SIGNAL n934 : STD_LOGIC;
   SIGNAL n935 : STD_LOGIC;
   SIGNAL n936 : STD_LOGIC;
   SIGNAL n937 : STD_LOGIC;
   SIGNAL n938 : STD_LOGIC;
   SIGNAL n939 : STD_LOGIC;
   SIGNAL n940 : STD_LOGIC;
   SIGNAL n1519 : STD_LOGIC;
   SIGNAL n1520 : STD_LOGIC;
   SIGNAL n1521 : STD_LOGIC;
   SIGNAL n1522 : STD_LOGIC;
   SIGNAL n1523 : STD_LOGIC;
   SIGNAL n1524 : STD_LOGIC;
   SIGNAL n1525 : STD_LOGIC;
   SIGNAL n1526 : STD_LOGIC;
   SIGNAL n1527 : STD_LOGIC;
   SIGNAL n1528 : STD_LOGIC;
   SIGNAL n1529 : STD_LOGIC;
   SIGNAL n1530 : STD_LOGIC;
   SIGNAL n1531 : STD_LOGIC;
   SIGNAL n1532 : STD_LOGIC;
   SIGNAL n1533 : STD_LOGIC;
   SIGNAL n1534 : STD_LOGIC;
   SIGNAL n1535 : STD_LOGIC;
   SIGNAL n1536 : STD_LOGIC;
   SIGNAL n1537 : STD_LOGIC;
   SIGNAL n1538 : STD_LOGIC;
   SIGNAL n1539 : STD_LOGIC;
   SIGNAL n1540 : STD_LOGIC;
   SIGNAL n1541 : STD_LOGIC;
   SIGNAL n1542 : STD_LOGIC;
   SIGNAL n1544 : STD_LOGIC;
   SIGNAL n1547 : STD_LOGIC;
   SIGNAL n1553 : STD_LOGIC;
   SIGNAL n1555 : STD_LOGIC;
   SIGNAL n2162 : STD_LOGIC;
   SIGNAL n2163 : STD_LOGIC;
   SIGNAL n2164 : STD_LOGIC;
   SIGNAL n2165 : STD_LOGIC;
   SIGNAL n2166 : STD_LOGIC;
   SIGNAL n2167 : STD_LOGIC;
   SIGNAL n2168 : STD_LOGIC;
   SIGNAL n2169 : STD_LOGIC;
   SIGNAL n2170 : STD_LOGIC;
   SIGNAL n2171 : STD_LOGIC;
   SIGNAL n2172 : STD_LOGIC;
   SIGNAL n2173 : STD_LOGIC;
   SIGNAL n2174 : STD_LOGIC;
   SIGNAL n2175 : STD_LOGIC;
   SIGNAL n2176 : STD_LOGIC;
   SIGNAL n2177 : STD_LOGIC;
   SIGNAL n2178 : STD_LOGIC;
   SIGNAL n2179 : STD_LOGIC;
   SIGNAL n2180 : STD_LOGIC;
   SIGNAL n2181 : STD_LOGIC;
   SIGNAL n2182 : STD_LOGIC;
   SIGNAL n2183 : STD_LOGIC;
   SIGNAL n2184 : STD_LOGIC;
   SIGNAL n2185 : STD_LOGIC;
   SIGNAL n2187 : STD_LOGIC;
   SIGNAL n2190 : STD_LOGIC;
   SIGNAL n2196 : STD_LOGIC;
   SIGNAL n2198 : STD_LOGIC;
   SIGNAL n2605 : STD_LOGIC;
   SIGNAL n2606 : STD_LOGIC;
   SIGNAL n2607 : STD_LOGIC;
   SIGNAL n2608 : STD_LOGIC;
   SIGNAL n2609 : STD_LOGIC;
   SIGNAL n2610 : STD_LOGIC;
   SIGNAL n2611 : STD_LOGIC;
   SIGNAL n2612 : STD_LOGIC;
   SIGNAL n2613 : STD_LOGIC;
   SIGNAL n2614 : STD_LOGIC;
   SIGNAL n2615 : STD_LOGIC;
   SIGNAL n2616 : STD_LOGIC;
   SIGNAL n2617 : STD_LOGIC;
   SIGNAL n2618 : STD_LOGIC;
   SIGNAL n2619 : STD_LOGIC;
   SIGNAL n2620 : STD_LOGIC;
   SIGNAL n2621 : STD_LOGIC;
   SIGNAL n2622 : STD_LOGIC;
   SIGNAL n2623 : STD_LOGIC;
   SIGNAL n2624 : STD_LOGIC;
   SIGNAL n2625 : STD_LOGIC;
   SIGNAL n2626 : STD_LOGIC;
   SIGNAL n2627 : STD_LOGIC;
   SIGNAL n2628 : STD_LOGIC;
   SIGNAL n2629 : STD_LOGIC;
   SIGNAL n2630 : STD_LOGIC;
   SIGNAL n2631 : STD_LOGIC;
   SIGNAL n2632 : STD_LOGIC;
   SIGNAL n2633 : STD_LOGIC;
   SIGNAL n2634 : STD_LOGIC;
   SIGNAL n2635 : STD_LOGIC;
   SIGNAL n2636 : STD_LOGIC;
   SIGNAL n2637 : STD_LOGIC;
   SIGNAL n2638 : STD_LOGIC;
   SIGNAL n2639 : STD_LOGIC;
   SIGNAL n2640 : STD_LOGIC;
   SIGNAL n2641 : STD_LOGIC;
   SIGNAL n2642 : STD_LOGIC;
   SIGNAL n2643 : STD_LOGIC;
   SIGNAL n2644 : STD_LOGIC;
   SIGNAL n2645 : STD_LOGIC;
   SIGNAL n2646 : STD_LOGIC;
   SIGNAL n2647 : STD_LOGIC;
   SIGNAL n2648 : STD_LOGIC;
   SIGNAL n2649 : STD_LOGIC;
   SIGNAL n2650 : STD_LOGIC;
   SIGNAL n2651 : STD_LOGIC;
   SIGNAL n2652 : STD_LOGIC;
   SIGNAL n2653 : STD_LOGIC;
   SIGNAL n2654 : STD_LOGIC;
   SIGNAL n2655 : STD_LOGIC;
   SIGNAL n2656 : STD_LOGIC;
   SIGNAL n2657 : STD_LOGIC;
   SIGNAL n2658 : STD_LOGIC;
   SIGNAL n2659 : STD_LOGIC;
   SIGNAL n2660 : STD_LOGIC;
   SIGNAL n2661 : STD_LOGIC;
   SIGNAL n2662 : STD_LOGIC;
   SIGNAL n2663 : STD_LOGIC;
   SIGNAL n2664 : STD_LOGIC;
   SIGNAL n2665 : STD_LOGIC;
   SIGNAL n2666 : STD_LOGIC;
   SIGNAL n2667 : STD_LOGIC;
   SIGNAL n2668 : STD_LOGIC;
   SIGNAL n2669 : STD_LOGIC;
   SIGNAL n2670 : STD_LOGIC;
   SIGNAL n2671 : STD_LOGIC;
   SIGNAL n2672 : STD_LOGIC;
   SIGNAL n2673 : STD_LOGIC;
   SIGNAL n2674 : STD_LOGIC;
   SIGNAL n2675 : STD_LOGIC;
   SIGNAL n2676 : STD_LOGIC;
   SIGNAL n2677 : STD_LOGIC;
   SIGNAL n2678 : STD_LOGIC;
   SIGNAL n2679 : STD_LOGIC;
   SIGNAL n2680 : STD_LOGIC;
   SIGNAL n2681 : STD_LOGIC;
   SIGNAL n2682 : STD_LOGIC;
   SIGNAL n2683 : STD_LOGIC;
   SIGNAL n2684 : STD_LOGIC;
   SIGNAL n2685 : STD_LOGIC;
   SIGNAL n2686 : STD_LOGIC;
   SIGNAL n2687 : STD_LOGIC;
   SIGNAL n2688 : STD_LOGIC;
   SIGNAL n2689 : STD_LOGIC;
   SIGNAL n2690 : STD_LOGIC;
   SIGNAL n2691 : STD_LOGIC;
   SIGNAL n2692 : STD_LOGIC;
   SIGNAL n2693 : STD_LOGIC;
   SIGNAL n2694 : STD_LOGIC;
   SIGNAL n2695 : STD_LOGIC;
   SIGNAL n2696 : STD_LOGIC;
   SIGNAL n2697 : STD_LOGIC;
   SIGNAL n2698 : STD_LOGIC;
   SIGNAL n2699 : STD_LOGIC;
   SIGNAL n2700 : STD_LOGIC;
   SIGNAL n2701 : STD_LOGIC;
   SIGNAL n2702 : STD_LOGIC;
   SIGNAL n2703 : STD_LOGIC;
   SIGNAL n2704 : STD_LOGIC;
   SIGNAL n2705 : STD_LOGIC;
   SIGNAL n2706 : STD_LOGIC;
   SIGNAL n2707 : STD_LOGIC;
   SIGNAL n2708 : STD_LOGIC;
   SIGNAL n2709 : STD_LOGIC;
   SIGNAL n2710 : STD_LOGIC;
   SIGNAL n2711 : STD_LOGIC;
   SIGNAL n2712 : STD_LOGIC;
   SIGNAL n2713 : STD_LOGIC;
   SIGNAL n2714 : STD_LOGIC;
   SIGNAL n2715 : STD_LOGIC;
   SIGNAL n2716 : STD_LOGIC;
   SIGNAL n2717 : STD_LOGIC;
   SIGNAL n2718 : STD_LOGIC;
   SIGNAL n2719 : STD_LOGIC;
   SIGNAL n2720 : STD_LOGIC;
   SIGNAL n2721 : STD_LOGIC;
   SIGNAL n2722 : STD_LOGIC;
   SIGNAL n2723 : STD_LOGIC;
   SIGNAL n2724 : STD_LOGIC;
   SIGNAL n2725 : STD_LOGIC;
   SIGNAL n2726 : STD_LOGIC;
   SIGNAL n2727 : STD_LOGIC;
   SIGNAL n2728 : STD_LOGIC;
   SIGNAL n2729 : STD_LOGIC;
   SIGNAL n2730 : STD_LOGIC;
   SIGNAL n2731 : STD_LOGIC;
   SIGNAL n2732 : STD_LOGIC;
   SIGNAL n2733 : STD_LOGIC;
   SIGNAL n2734 : STD_LOGIC;
   SIGNAL n2735 : STD_LOGIC;
   SIGNAL n2736 : STD_LOGIC;
   SIGNAL n2737 : STD_LOGIC;
   SIGNAL n2738 : STD_LOGIC;
   SIGNAL n2739 : STD_LOGIC;
   SIGNAL n2740 : STD_LOGIC;
   SIGNAL n2741 : STD_LOGIC;
   SIGNAL n2742 : STD_LOGIC;
   SIGNAL n2743 : STD_LOGIC;
   SIGNAL n2744 : STD_LOGIC;
   SIGNAL n2745 : STD_LOGIC;
   SIGNAL n2746 : STD_LOGIC;
   SIGNAL n2747 : STD_LOGIC;
   SIGNAL n2748 : STD_LOGIC;
   SIGNAL n2749 : STD_LOGIC;
   SIGNAL n2750 : STD_LOGIC;
   SIGNAL n2751 : STD_LOGIC;
   SIGNAL n2752 : STD_LOGIC;
   SIGNAL n2753 : STD_LOGIC;
   SIGNAL n2754 : STD_LOGIC;
   SIGNAL n2755 : STD_LOGIC;
   SIGNAL n2756 : STD_LOGIC;
   SIGNAL n2757 : STD_LOGIC;
   SIGNAL n2758 : STD_LOGIC;
   SIGNAL n2759 : STD_LOGIC;
   SIGNAL n2760 : STD_LOGIC;
   SIGNAL n2761 : STD_LOGIC;
   SIGNAL n2762 : STD_LOGIC;
   SIGNAL n2763 : STD_LOGIC;
   SIGNAL n2764 : STD_LOGIC;
   SIGNAL n2765 : STD_LOGIC;
   SIGNAL n2766 : STD_LOGIC;
   SIGNAL n2767 : STD_LOGIC;
   SIGNAL n2768 : STD_LOGIC;
   SIGNAL n2769 : STD_LOGIC;
   SIGNAL n2770 : STD_LOGIC;
   SIGNAL n2771 : STD_LOGIC;
   SIGNAL n2772 : STD_LOGIC;
   SIGNAL n2773 : STD_LOGIC;
   SIGNAL n3014 : STD_LOGIC;
   SIGNAL n3015 : STD_LOGIC;
   SIGNAL n3016 : STD_LOGIC;
   SIGNAL n3017 : STD_LOGIC;
   SIGNAL n3018 : STD_LOGIC;
   SIGNAL n3019 : STD_LOGIC;
   SIGNAL n3020 : STD_LOGIC;
   SIGNAL n3021 : STD_LOGIC;
   SIGNAL n3022 : STD_LOGIC;
   SIGNAL n3023 : STD_LOGIC;
   SIGNAL n3024 : STD_LOGIC;
   SIGNAL n3025 : STD_LOGIC;
   SIGNAL n3026 : STD_LOGIC;
   SIGNAL n3027 : STD_LOGIC;
   SIGNAL n3028 : STD_LOGIC;
   SIGNAL n3029 : STD_LOGIC;
   SIGNAL n3030 : STD_LOGIC;
   SIGNAL n3031 : STD_LOGIC;
   SIGNAL n3032 : STD_LOGIC;
   SIGNAL n3033 : STD_LOGIC;
   SIGNAL n3034 : STD_LOGIC;
   SIGNAL n3035 : STD_LOGIC;
   SIGNAL n3036 : STD_LOGIC;
   SIGNAL n3037 : STD_LOGIC;
   SIGNAL n3039 : STD_LOGIC;
   SIGNAL n3042 : STD_LOGIC;
   SIGNAL n3066 : STD_LOGIC;
   SIGNAL n3068 : STD_LOGIC;
   SIGNAL n3531 : STD_LOGIC;
   SIGNAL n3532 : STD_LOGIC;
   SIGNAL n3533 : STD_LOGIC;
   SIGNAL n3534 : STD_LOGIC;
   SIGNAL n3535 : STD_LOGIC;
   SIGNAL n3536 : STD_LOGIC;
   SIGNAL n3537 : STD_LOGIC;
   SIGNAL n3538 : STD_LOGIC;
   SIGNAL n3539 : STD_LOGIC;
   SIGNAL n3540 : STD_LOGIC;
   SIGNAL n3541 : STD_LOGIC;
   SIGNAL n3542 : STD_LOGIC;
   SIGNAL n3543 : STD_LOGIC;
   SIGNAL n3544 : STD_LOGIC;
   SIGNAL n3545 : STD_LOGIC;
   SIGNAL n3546 : STD_LOGIC;
   SIGNAL n3547 : STD_LOGIC;
   SIGNAL n3548 : STD_LOGIC;
   SIGNAL n3549 : STD_LOGIC;
   SIGNAL n3550 : STD_LOGIC;
   SIGNAL n3551 : STD_LOGIC;
   SIGNAL n3552 : STD_LOGIC;
   SIGNAL n3553 : STD_LOGIC;
   SIGNAL n3554 : STD_LOGIC;
   SIGNAL n3556 : STD_LOGIC;
   SIGNAL n3559 : STD_LOGIC;
   SIGNAL n3583 : STD_LOGIC;
   SIGNAL n3585 : STD_LOGIC;
   SIGNAL n4445 : STD_LOGIC;
   SIGNAL n6691 : STD_LOGIC;
   SIGNAL n6692 : STD_LOGIC;
   SIGNAL n6693 : STD_LOGIC;
   SIGNAL n6694 : STD_LOGIC;
   SIGNAL n6695 : STD_LOGIC;
   SIGNAL n6696 : STD_LOGIC;
   SIGNAL n6697 : STD_LOGIC;
   SIGNAL n6698 : STD_LOGIC;
   SIGNAL n6699 : STD_LOGIC;
   SIGNAL n6700 : STD_LOGIC;
   SIGNAL n6701 : STD_LOGIC;
   SIGNAL n6702 : STD_LOGIC;
   SIGNAL n6703 : STD_LOGIC;
   SIGNAL n6704 : STD_LOGIC;
   SIGNAL n6705 : STD_LOGIC;
   SIGNAL n6706 : STD_LOGIC;
   SIGNAL n6707 : STD_LOGIC;
   SIGNAL n6708 : STD_LOGIC;
   SIGNAL n6709 : STD_LOGIC;
   SIGNAL n6710 : STD_LOGIC;
   SIGNAL n6711 : STD_LOGIC;
   SIGNAL n6712 : STD_LOGIC;
   SIGNAL n6713 : STD_LOGIC;
   SIGNAL n6714 : STD_LOGIC;
   SIGNAL n6715 : STD_LOGIC;
   SIGNAL n6716 : STD_LOGIC;
   SIGNAL n6717 : STD_LOGIC;
   SIGNAL n6718 : STD_LOGIC;
   SIGNAL n6719 : STD_LOGIC;
   SIGNAL n6720 : STD_LOGIC;
   SIGNAL n6721 : STD_LOGIC;
   SIGNAL n6722 : STD_LOGIC;
   SIGNAL n6723 : STD_LOGIC;
   SIGNAL n6724 : STD_LOGIC;
   SIGNAL n6725 : STD_LOGIC;
   SIGNAL n6726 : STD_LOGIC;
   SIGNAL n6727 : STD_LOGIC;
   SIGNAL n6728 : STD_LOGIC;
   SIGNAL n6729 : STD_LOGIC;
   SIGNAL n6730 : STD_LOGIC;
   SIGNAL n6731 : STD_LOGIC;
   SIGNAL n6732 : STD_LOGIC;
   SIGNAL n6733 : STD_LOGIC;
   SIGNAL n6734 : STD_LOGIC;
   SIGNAL n6735 : STD_LOGIC;
   SIGNAL n6736 : STD_LOGIC;
   SIGNAL n6737 : STD_LOGIC;
   SIGNAL n6738 : STD_LOGIC;
   SIGNAL n6739 : STD_LOGIC;
   SIGNAL n6740 : STD_LOGIC;
   SIGNAL n6741 : STD_LOGIC;
   SIGNAL n6742 : STD_LOGIC;
   SIGNAL n6743 : STD_LOGIC;
   SIGNAL n6744 : STD_LOGIC;
   SIGNAL n6745 : STD_LOGIC;
   SIGNAL n6746 : STD_LOGIC;
   SIGNAL n6747 : STD_LOGIC;
   SIGNAL n6748 : STD_LOGIC;
   SIGNAL n6749 : STD_LOGIC;
   SIGNAL n6750 : STD_LOGIC;
   SIGNAL n6751 : STD_LOGIC;
   SIGNAL n6752 : STD_LOGIC;
   SIGNAL n6753 : STD_LOGIC;
   SIGNAL n6754 : STD_LOGIC;
   SIGNAL n6755 : STD_LOGIC;
   SIGNAL n6756 : STD_LOGIC;
   SIGNAL n6757 : STD_LOGIC;
   SIGNAL n6758 : STD_LOGIC;
   SIGNAL n6759 : STD_LOGIC;
   SIGNAL n6760 : STD_LOGIC;
   SIGNAL n6761 : STD_LOGIC;
   SIGNAL n6762 : STD_LOGIC;
   SIGNAL n6763 : STD_LOGIC;
   SIGNAL n6815 : STD_LOGIC;
   SIGNAL n6816 : STD_LOGIC;
   SIGNAL n6817 : STD_LOGIC;
   SIGNAL n6818 : STD_LOGIC;
   SIGNAL n6819 : STD_LOGIC;
   SIGNAL n6820 : STD_LOGIC;
   SIGNAL n6821 : STD_LOGIC;
   SIGNAL n7164 : STD_LOGIC;
   SIGNAL n7277 : STD_LOGIC;
   SIGNAL n7278 : STD_LOGIC;
   SIGNAL n7279 : STD_LOGIC;
   SIGNAL n7280 : STD_LOGIC;
   SIGNAL n7281 : STD_LOGIC;
   SIGNAL n7282 : STD_LOGIC;
   SIGNAL n7283 : STD_LOGIC;
   SIGNAL n7284 : STD_LOGIC;
   SIGNAL n7285 : STD_LOGIC;
   SIGNAL n7286 : STD_LOGIC;
   SIGNAL n7287 : STD_LOGIC;
   SIGNAL n7288 : STD_LOGIC;
   SIGNAL n7289 : STD_LOGIC;
   SIGNAL n7290 : STD_LOGIC;
   SIGNAL n7291 : STD_LOGIC;
   SIGNAL n7292 : STD_LOGIC;
   SIGNAL n7294 : STD_LOGIC;
   SIGNAL n7297 : STD_LOGIC;
   SIGNAL n7325 : STD_LOGIC;
   SIGNAL n7327 : STD_LOGIC;
   SIGNAL n7834 : STD_LOGIC;
   SIGNAL n7835 : STD_LOGIC;
   SIGNAL n7836 : STD_LOGIC;
   SIGNAL n7837 : STD_LOGIC;
   SIGNAL n7838 : STD_LOGIC;
   SIGNAL n7839 : STD_LOGIC;
   SIGNAL n7840 : STD_LOGIC;
   SIGNAL n7841 : STD_LOGIC;
   SIGNAL n7842 : STD_LOGIC;
   SIGNAL n7843 : STD_LOGIC;
   SIGNAL n7844 : STD_LOGIC;
   SIGNAL n7845 : STD_LOGIC;
   SIGNAL n7846 : STD_LOGIC;
   SIGNAL n7847 : STD_LOGIC;
   SIGNAL n7848 : STD_LOGIC;
   SIGNAL n7849 : STD_LOGIC;
   SIGNAL n7850 : STD_LOGIC;
   SIGNAL n7851 : STD_LOGIC;
   SIGNAL n7852 : STD_LOGIC;
   SIGNAL n7853 : STD_LOGIC;
   SIGNAL n7854 : STD_LOGIC;
   SIGNAL n7855 : STD_LOGIC;
   SIGNAL n7856 : STD_LOGIC;
   SIGNAL n7857 : STD_LOGIC;
   SIGNAL n7858 : STD_LOGIC;
   SIGNAL n7859 : STD_LOGIC;
   SIGNAL n7860 : STD_LOGIC;
   SIGNAL n7861 : STD_LOGIC;
   SIGNAL n7862 : STD_LOGIC;
   SIGNAL n7863 : STD_LOGIC;
   SIGNAL n7865 : STD_LOGIC;
   SIGNAL n7868 : STD_LOGIC;
   SIGNAL n7874 : STD_LOGIC;
   SIGNAL n7876 : STD_LOGIC;
   SIGNAL n8379 : STD_LOGIC;
   SIGNAL n8380 : STD_LOGIC;
   SIGNAL n8381 : STD_LOGIC;
   SIGNAL n8382 : STD_LOGIC;
   SIGNAL n8383 : STD_LOGIC;
   SIGNAL n8384 : STD_LOGIC;
   SIGNAL n8385 : STD_LOGIC;
   SIGNAL n8386 : STD_LOGIC;
   SIGNAL n8387 : STD_LOGIC;
   SIGNAL n8388 : STD_LOGIC;
   SIGNAL n8389 : STD_LOGIC;
   SIGNAL n8390 : STD_LOGIC;
   SIGNAL n8391 : STD_LOGIC;
   SIGNAL n8392 : STD_LOGIC;
   SIGNAL n8393 : STD_LOGIC;
   SIGNAL n8394 : STD_LOGIC;
   SIGNAL n8395 : STD_LOGIC;
   SIGNAL n8396 : STD_LOGIC;
   SIGNAL n8397 : STD_LOGIC;
   SIGNAL n8398 : STD_LOGIC;
   SIGNAL n8399 : STD_LOGIC;
   SIGNAL n8400 : STD_LOGIC;
   SIGNAL n8401 : STD_LOGIC;
   SIGNAL n8402 : STD_LOGIC;
   SIGNAL n8403 : STD_LOGIC;
   SIGNAL n8404 : STD_LOGIC;
   SIGNAL n8405 : STD_LOGIC;
   SIGNAL n8406 : STD_LOGIC;
   SIGNAL n8407 : STD_LOGIC;
   SIGNAL n8408 : STD_LOGIC;
   SIGNAL n8410 : STD_LOGIC;
   SIGNAL n8413 : STD_LOGIC;
   SIGNAL n8419 : STD_LOGIC;
   SIGNAL n8421 : STD_LOGIC;

BEGIN

   n138 <= DIN(0);
   n139 <= DIN(1);
   n140 <= DIN(2);
   n141 <= DIN(3);
   n142 <= DIN(4);
   n143 <= DIN(5);
   n144 <= DIN(6);
   n145 <= DIN(7);
   n146 <= DIN(8);
   n147 <= DIN(9);
   n148 <= DIN(10);
   n149 <= DIN(11);
   n150 <= DIN(12);
   n151 <= DIN(13);
   n152 <= ND;
   n155 <= CLK;
   n156 <= ADDR(0);
   n157 <= ADDR(1);
   n158 <= ADDR(2);
   n159 <= ADDR(3);
   n160 <= ADDR(4);
   n161 <= LD_DIN(0);
   n162 <= LD_DIN(1);
   n163 <= LD_DIN(2);
   n164 <= LD_DIN(3);
   n165 <= LD_DIN(4);
   n166 <= LD_DIN(5);
   n167 <= LD_DIN(6);
   n168 <= LD_DIN(7);
   n169 <= LD_DIN(8);
   n170 <= LD_DIN(9);
   n171 <= LD_DIN(10);
   n172 <= LD_DIN(11);
   n173 <= LD_DIN(12);
   n174 <= LD_DIN(13);
   n175 <= LD_DIN(14);
   n176 <= LD_DIN(15);
   n177 <= LD_DIN(16);
   n178 <= LD_DIN(17);
   n179 <= LD_DIN(18);
   n180 <= LD_DIN(19);
   n181 <= LD_DIN(20);
   n182 <= LD_DIN(21);
   n183 <= LD_DIN(22);
   n184 <= LD_DIN(23);
   n185 <= LD_DIN(24);
   n186 <= LD_DIN(25);
   n187 <= LD_DIN(26);
   n188 <= LD_DIN(27);
   n189 <= LD_DIN(28);
   n190 <= LD_DIN(29);
   n191 <= LD_DIN(30);
   n192 <= LD_DIN(31);
   n193 <= WE;
   n194 <= SEL;
   RDY <= n153;
   RFD <= n154;
   DOUT_I(0) <= n195;
   DOUT_I(1) <= n196;
   DOUT_I(2) <= n197;
   DOUT_I(3) <= n198;
   DOUT_I(4) <= n199;
   DOUT_I(5) <= n200;
   DOUT_I(6) <= n201;
   DOUT_I(7) <= n202;
   DOUT_I(8) <= n203;
   DOUT_I(9) <= n204;
   DOUT_I(10) <= n205;
   DOUT_I(11) <= n206;
   DOUT_I(12) <= n207;
   DOUT_I(13) <= n208;
   DOUT_I(14) <= n209;
   DOUT_I(15) <= n210;
   DOUT_I(16) <= n211;
   DOUT_I(17) <= n212;
   DOUT_I(18) <= n213;
   DOUT_I(19) <= n214;
   DOUT_I(20) <= n215;
   DOUT_I(21) <= n216;
   DOUT_I(22) <= n217;
   DOUT_I(23) <= n218;
   DOUT_I(24) <= n219;
   DOUT_I(25) <= n220;
   DOUT_I(26) <= n221;
   DOUT_I(27) <= n222;
   DOUT_I(28) <= n223;
   DOUT_I(29) <= n224;
   DOUT_Q(0) <= n225;
   DOUT_Q(1) <= n226;
   DOUT_Q(2) <= n227;
   DOUT_Q(3) <= n228;
   DOUT_Q(4) <= n229;
   DOUT_Q(5) <= n230;
   DOUT_Q(6) <= n231;
   DOUT_Q(7) <= n232;
   DOUT_Q(8) <= n233;
   DOUT_Q(9) <= n234;
   DOUT_Q(10) <= n235;
   DOUT_Q(11) <= n236;
   DOUT_Q(12) <= n237;
   DOUT_Q(13) <= n238;
   DOUT_Q(14) <= n239;
   DOUT_Q(15) <= n240;
   DOUT_Q(16) <= n241;
   DOUT_Q(17) <= n242;
   DOUT_Q(18) <= n243;
   DOUT_Q(19) <= n244;
   DOUT_Q(20) <= n245;
   DOUT_Q(21) <= n246;
   DOUT_Q(22) <= n247;
   DOUT_Q(23) <= n248;
   DOUT_Q(24) <= n249;
   DOUT_Q(25) <= n250;
   DOUT_Q(26) <= n251;
   DOUT_Q(27) <= n252;
   DOUT_Q(28) <= n253;
   DOUT_Q(29) <= n254;

   BU4_I0 <= n160;
   BU4_I1 <= n159;
   BU4_I2 <= n158;
   BU4_I3 <= n194;
   n54 <= BU4_O;
   BU4 : LUT4
      GENERIC MAP (
         INIT  => X"1000"
      )
      PORT MAP (
         I0 => BU4_I0,
         I1 => BU4_I1,
         I2 => BU4_I2,
         I3 => BU4_I3,
         O => BU4_O
      );

   BU8_I0 <= n54;
   BU8_I1 <= n193;
   BU8_I2 <= n157;
   BU8_I3 <= n156;
   n294 <= BU8_O;
   BU8 : LUT4
      GENERIC MAP (
         INIT  => X"0080"
      )
      PORT MAP (
         I0 => BU8_I0,
         I1 => BU8_I1,
         I2 => BU8_I2,
         I3 => BU8_I3,
         O => BU8_O
      );

   BU10_I0 <= '1';
   BU10_I1 <= '0';
   BU10_I2 <= '0';
   BU10_I3 <= '0';
   n154 <= BU10_O;
   BU10 : LUT4
      GENERIC MAP (
         INIT  => X"aaaa"
      )
      PORT MAP (
         I0 => BU10_I0,
         I1 => BU10_I1,
         I2 => BU10_I2,
         I3 => BU10_I3,
         O => BU10_O
      );

   BU1292_D <= n152;
   BU1292_C <= n155;
   BU1292_CE <= '1';
   n343 <= BU1292_Q;
   BU1292 : FDE
      PORT MAP (
         D => BU1292_D,
         C => BU1292_C,
         CE => BU1292_CE,
         Q => BU1292_Q
      );

   BU14_D <= n138;
   BU14_CE <= n152;
   BU14_CLK <= n155;
   BU14_A0 <= '0';
   BU14_A1 <= '1';
   BU14_A2 <= '0';
   BU14_A3 <= '0';
   n927 <= BU14_Q;
   BU14 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU14_D,
         CE => BU14_CE,
         CLK => BU14_CLK,
         A0 => BU14_A0,
         A1 => BU14_A1,
         A2 => BU14_A2,
         A3 => BU14_A3,
         Q => BU14_Q
      );

   BU16_D <= n927;
   BU16_C <= n155;
   BU16_CE <= n152;
   n590 <= BU16_Q;
   BU16 : FDE
      PORT MAP (
         D => BU16_D,
         C => BU16_C,
         CE => BU16_CE,
         Q => BU16_Q
      );

   BU17_D <= n139;
   BU17_CE <= n152;
   BU17_CLK <= n155;
   BU17_A0 <= '0';
   BU17_A1 <= '1';
   BU17_A2 <= '0';
   BU17_A3 <= '0';
   n928 <= BU17_Q;
   BU17 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU17_D,
         CE => BU17_CE,
         CLK => BU17_CLK,
         A0 => BU17_A0,
         A1 => BU17_A1,
         A2 => BU17_A2,
         A3 => BU17_A3,
         Q => BU17_Q
      );

   BU19_D <= n928;
   BU19_C <= n155;
   BU19_CE <= n152;
   n589 <= BU19_Q;
   BU19 : FDE
      PORT MAP (
         D => BU19_D,
         C => BU19_C,
         CE => BU19_CE,
         Q => BU19_Q
      );

   BU20_D <= n140;
   BU20_CE <= n152;
   BU20_CLK <= n155;
   BU20_A0 <= '0';
   BU20_A1 <= '1';
   BU20_A2 <= '0';
   BU20_A3 <= '0';
   n929 <= BU20_Q;
   BU20 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU20_D,
         CE => BU20_CE,
         CLK => BU20_CLK,
         A0 => BU20_A0,
         A1 => BU20_A1,
         A2 => BU20_A2,
         A3 => BU20_A3,
         Q => BU20_Q
      );

   BU22_D <= n929;
   BU22_C <= n155;
   BU22_CE <= n152;
   n588 <= BU22_Q;
   BU22 : FDE
      PORT MAP (
         D => BU22_D,
         C => BU22_C,
         CE => BU22_CE,
         Q => BU22_Q
      );

   BU23_D <= n141;
   BU23_CE <= n152;
   BU23_CLK <= n155;
   BU23_A0 <= '0';
   BU23_A1 <= '1';
   BU23_A2 <= '0';
   BU23_A3 <= '0';
   n930 <= BU23_Q;
   BU23 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU23_D,
         CE => BU23_CE,
         CLK => BU23_CLK,
         A0 => BU23_A0,
         A1 => BU23_A1,
         A2 => BU23_A2,
         A3 => BU23_A3,
         Q => BU23_Q
      );

   BU25_D <= n930;
   BU25_C <= n155;
   BU25_CE <= n152;
   n587 <= BU25_Q;
   BU25 : FDE
      PORT MAP (
         D => BU25_D,
         C => BU25_C,
         CE => BU25_CE,
         Q => BU25_Q
      );

   BU26_D <= n142;
   BU26_CE <= n152;
   BU26_CLK <= n155;
   BU26_A0 <= '0';
   BU26_A1 <= '1';
   BU26_A2 <= '0';
   BU26_A3 <= '0';
   n931 <= BU26_Q;
   BU26 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU26_D,
         CE => BU26_CE,
         CLK => BU26_CLK,
         A0 => BU26_A0,
         A1 => BU26_A1,
         A2 => BU26_A2,
         A3 => BU26_A3,
         Q => BU26_Q
      );

   BU28_D <= n931;
   BU28_C <= n155;
   BU28_CE <= n152;
   n586 <= BU28_Q;
   BU28 : FDE
      PORT MAP (
         D => BU28_D,
         C => BU28_C,
         CE => BU28_CE,
         Q => BU28_Q
      );

   BU29_D <= n143;
   BU29_CE <= n152;
   BU29_CLK <= n155;
   BU29_A0 <= '0';
   BU29_A1 <= '1';
   BU29_A2 <= '0';
   BU29_A3 <= '0';
   n932 <= BU29_Q;
   BU29 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU29_D,
         CE => BU29_CE,
         CLK => BU29_CLK,
         A0 => BU29_A0,
         A1 => BU29_A1,
         A2 => BU29_A2,
         A3 => BU29_A3,
         Q => BU29_Q
      );

   BU31_D <= n932;
   BU31_C <= n155;
   BU31_CE <= n152;
   n585 <= BU31_Q;
   BU31 : FDE
      PORT MAP (
         D => BU31_D,
         C => BU31_C,
         CE => BU31_CE,
         Q => BU31_Q
      );

   BU32_D <= n144;
   BU32_CE <= n152;
   BU32_CLK <= n155;
   BU32_A0 <= '0';
   BU32_A1 <= '1';
   BU32_A2 <= '0';
   BU32_A3 <= '0';
   n933 <= BU32_Q;
   BU32 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU32_D,
         CE => BU32_CE,
         CLK => BU32_CLK,
         A0 => BU32_A0,
         A1 => BU32_A1,
         A2 => BU32_A2,
         A3 => BU32_A3,
         Q => BU32_Q
      );

   BU34_D <= n933;
   BU34_C <= n155;
   BU34_CE <= n152;
   n584 <= BU34_Q;
   BU34 : FDE
      PORT MAP (
         D => BU34_D,
         C => BU34_C,
         CE => BU34_CE,
         Q => BU34_Q
      );

   BU35_D <= n145;
   BU35_CE <= n152;
   BU35_CLK <= n155;
   BU35_A0 <= '0';
   BU35_A1 <= '1';
   BU35_A2 <= '0';
   BU35_A3 <= '0';
   n934 <= BU35_Q;
   BU35 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU35_D,
         CE => BU35_CE,
         CLK => BU35_CLK,
         A0 => BU35_A0,
         A1 => BU35_A1,
         A2 => BU35_A2,
         A3 => BU35_A3,
         Q => BU35_Q
      );

   BU37_D <= n934;
   BU37_C <= n155;
   BU37_CE <= n152;
   n583 <= BU37_Q;
   BU37 : FDE
      PORT MAP (
         D => BU37_D,
         C => BU37_C,
         CE => BU37_CE,
         Q => BU37_Q
      );

   BU38_D <= n146;
   BU38_CE <= n152;
   BU38_CLK <= n155;
   BU38_A0 <= '0';
   BU38_A1 <= '1';
   BU38_A2 <= '0';
   BU38_A3 <= '0';
   n935 <= BU38_Q;
   BU38 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU38_D,
         CE => BU38_CE,
         CLK => BU38_CLK,
         A0 => BU38_A0,
         A1 => BU38_A1,
         A2 => BU38_A2,
         A3 => BU38_A3,
         Q => BU38_Q
      );

   BU40_D <= n935;
   BU40_C <= n155;
   BU40_CE <= n152;
   n582 <= BU40_Q;
   BU40 : FDE
      PORT MAP (
         D => BU40_D,
         C => BU40_C,
         CE => BU40_CE,
         Q => BU40_Q
      );

   BU41_D <= n147;
   BU41_CE <= n152;
   BU41_CLK <= n155;
   BU41_A0 <= '0';
   BU41_A1 <= '1';
   BU41_A2 <= '0';
   BU41_A3 <= '0';
   n936 <= BU41_Q;
   BU41 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU41_D,
         CE => BU41_CE,
         CLK => BU41_CLK,
         A0 => BU41_A0,
         A1 => BU41_A1,
         A2 => BU41_A2,
         A3 => BU41_A3,
         Q => BU41_Q
      );

   BU43_D <= n936;
   BU43_C <= n155;
   BU43_CE <= n152;
   n581 <= BU43_Q;
   BU43 : FDE
      PORT MAP (
         D => BU43_D,
         C => BU43_C,
         CE => BU43_CE,
         Q => BU43_Q
      );

   BU44_D <= n148;
   BU44_CE <= n152;
   BU44_CLK <= n155;
   BU44_A0 <= '0';
   BU44_A1 <= '1';
   BU44_A2 <= '0';
   BU44_A3 <= '0';
   n937 <= BU44_Q;
   BU44 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU44_D,
         CE => BU44_CE,
         CLK => BU44_CLK,
         A0 => BU44_A0,
         A1 => BU44_A1,
         A2 => BU44_A2,
         A3 => BU44_A3,
         Q => BU44_Q
      );

   BU46_D <= n937;
   BU46_C <= n155;
   BU46_CE <= n152;
   n580 <= BU46_Q;
   BU46 : FDE
      PORT MAP (
         D => BU46_D,
         C => BU46_C,
         CE => BU46_CE,
         Q => BU46_Q
      );

   BU47_D <= n149;
   BU47_CE <= n152;
   BU47_CLK <= n155;
   BU47_A0 <= '0';
   BU47_A1 <= '1';
   BU47_A2 <= '0';
   BU47_A3 <= '0';
   n938 <= BU47_Q;
   BU47 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU47_D,
         CE => BU47_CE,
         CLK => BU47_CLK,
         A0 => BU47_A0,
         A1 => BU47_A1,
         A2 => BU47_A2,
         A3 => BU47_A3,
         Q => BU47_Q
      );

   BU49_D <= n938;
   BU49_C <= n155;
   BU49_CE <= n152;
   n579 <= BU49_Q;
   BU49 : FDE
      PORT MAP (
         D => BU49_D,
         C => BU49_C,
         CE => BU49_CE,
         Q => BU49_Q
      );

   BU50_D <= n150;
   BU50_CE <= n152;
   BU50_CLK <= n155;
   BU50_A0 <= '0';
   BU50_A1 <= '1';
   BU50_A2 <= '0';
   BU50_A3 <= '0';
   n939 <= BU50_Q;
   BU50 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU50_D,
         CE => BU50_CE,
         CLK => BU50_CLK,
         A0 => BU50_A0,
         A1 => BU50_A1,
         A2 => BU50_A2,
         A3 => BU50_A3,
         Q => BU50_Q
      );

   BU52_D <= n939;
   BU52_C <= n155;
   BU52_CE <= n152;
   n578 <= BU52_Q;
   BU52 : FDE
      PORT MAP (
         D => BU52_D,
         C => BU52_C,
         CE => BU52_CE,
         Q => BU52_Q
      );

   BU53_D <= n151;
   BU53_CE <= n152;
   BU53_CLK <= n155;
   BU53_A0 <= '0';
   BU53_A1 <= '1';
   BU53_A2 <= '0';
   BU53_A3 <= '0';
   n940 <= BU53_Q;
   BU53 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU53_D,
         CE => BU53_CE,
         CLK => BU53_CLK,
         A0 => BU53_A0,
         A1 => BU53_A1,
         A2 => BU53_A2,
         A3 => BU53_A3,
         Q => BU53_Q
      );

   BU55_D <= n940;
   BU55_C <= n155;
   BU55_CE <= n152;
   n577 <= BU55_Q;
   BU55 : FDE
      PORT MAP (
         D => BU55_D,
         C => BU55_C,
         CE => BU55_CE,
         Q => BU55_Q
      );

   BU57_DATA(0) <= n161;
   BU57_DATA(1) <= n162;
   BU57_DATA(2) <= n163;
   BU57_DATA(3) <= n164;
   BU57_DATA(4) <= n165;
   BU57_DATA(5) <= n166;
   BU57_DATA(6) <= n167;
   BU57_DATA(7) <= n168;
   BU57_DATA(8) <= n169;
   BU57_DATA(9) <= n170;
   BU57_DATA(10) <= n171;
   BU57_DATA(11) <= n172;
   BU57_DATA(12) <= n173;
   BU57_DATA(13) <= n174;
   BU57_DATA(14) <= n175;
   BU57_DATA(15) <= n176;
   BU57_DATA(16) <= n177;
   BU57_DATA(17) <= n178;
   BU57_DATA(18) <= n179;
   BU57_DATA(19) <= n180;
   BU57_DATA(20) <= n181;
   BU57_DATA(21) <= n182;
   BU57_DATA(22) <= n183;
   BU57_DATA(23) <= n184;
   BU57_DATA(24) <= n185;
   BU57_DATA(25) <= n186;
   BU57_DATA(26) <= n187;
   BU57_DATA(27) <= n188;
   BU57_DATA(28) <= n189;
   BU57_DATA(29) <= n190;
   BU57_DATA(30) <= n191;
   BU57_DATA(31) <= n192;
   BU57_WE <= n294;
   BU57_CLK <= n155;
   BU57_CE <= n152;
   n342 <= BU57_RDY;
   n429 <= BU57_SINE(0);
   n428 <= BU57_SINE(1);
   n427 <= BU57_SINE(2);
   n426 <= BU57_SINE(3);
   n425 <= BU57_SINE(4);
   n424 <= BU57_SINE(5);
   n423 <= BU57_SINE(6);
   n422 <= BU57_SINE(7);
   n421 <= BU57_SINE(8);
   n420 <= BU57_SINE(9);
   n419 <= BU57_SINE(10);
   n418 <= BU57_SINE(11);
   n417 <= BU57_SINE(12);
   n416 <= BU57_SINE(13);
   n415 <= BU57_SINE(14);
   n633 <= BU57_COSINE(0);
   n632 <= BU57_COSINE(1);
   n631 <= BU57_COSINE(2);
   n630 <= BU57_COSINE(3);
   n629 <= BU57_COSINE(4);
   n628 <= BU57_COSINE(5);
   n627 <= BU57_COSINE(6);
   n626 <= BU57_COSINE(7);
   n625 <= BU57_COSINE(8);
   n624 <= BU57_COSINE(9);
   n623 <= BU57_COSINE(10);
   n622 <= BU57_COSINE(11);
   n621 <= BU57_COSINE(12);
   n620 <= BU57_COSINE(13);
   n619 <= BU57_COSINE(14);
   BU57 : C_DDS_V4_1
      GENERIC MAP (
         c_phase_offset_value => "00000000000000000000000000000000",
         c_phase_increment_value => "01001100110011001100110011001101",
         c_has_rdy => 1,
         c_has_sclr => 0,
         c_phase_offset => 0,
         c_data_width => 32,
         c_accumulator_latency => 1,
         c_enable_rlocs => 0,
         c_phase_angle_width => 13,
         c_has_rfd => 0,
         c_phase_increment => 1,
         c_negative_sine => 0,
         c_latency => 4,
         c_has_ce => 1,
         c_has_aclr => 0,
         c_outputs_required => 2,
         c_pipelined => 1,
         c_accumulator_width => 32,
         c_mem_type => 1,
         c_negative_cosine => 0,
         c_noise_shaping => 1,
         c_output_width => 15
      )
      PORT MAP (
         DATA => BU57_DATA,
         WE => BU57_WE,
         CLK => BU57_CLK,
         CE => BU57_CE,
         RDY => BU57_RDY,
         SINE => BU57_SINE,
         COSINE => BU57_COSINE
      );

   BU1294_I0 <= n342;
   BU1294_I1 <= n343;
   BU1294_I2 <= '0';
   BU1294_I3 <= '0';
   n341 <= BU1294_O;
   BU1294 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU1294_I0,
         I1 => BU1294_I1,
         I2 => BU1294_I2,
         I3 => BU1294_I3,
         O => BU1294_O
      );

   BU1296_clk <= n155;
   BU1296_a(13) <= n577;
   BU1296_a(12) <= n578;
   BU1296_a(11) <= n579;
   BU1296_a(10) <= n580;
   BU1296_a(9) <= n581;
   BU1296_a(8) <= n582;
   BU1296_a(7) <= n583;
   BU1296_a(6) <= n584;
   BU1296_a(5) <= n585;
   BU1296_a(4) <= n586;
   BU1296_a(3) <= n587;
   BU1296_a(2) <= n588;
   BU1296_a(1) <= n589;
   BU1296_a(0) <= n590;
   BU1296_b(14) <= n415;
   BU1296_b(13) <= n416;
   BU1296_b(12) <= n417;
   BU1296_b(11) <= n418;
   BU1296_b(10) <= n419;
   BU1296_b(9) <= n420;
   BU1296_b(8) <= n421;
   BU1296_b(7) <= n422;
   BU1296_b(6) <= n423;
   BU1296_b(5) <= n424;
   BU1296_b(4) <= n425;
   BU1296_b(3) <= n426;
   BU1296_b(2) <= n427;
   BU1296_b(1) <= n428;
   BU1296_b(0) <= n429;
   n460 <= BU1296_q(28);
   n461 <= BU1296_q(27);
   n462 <= BU1296_q(26);
   n463 <= BU1296_q(25);
   n464 <= BU1296_q(24);
   n465 <= BU1296_q(23);
   n466 <= BU1296_q(22);
   n467 <= BU1296_q(21);
   n468 <= BU1296_q(20);
   n469 <= BU1296_q(19);
   n470 <= BU1296_q(18);
   n471 <= BU1296_q(17);
   n472 <= BU1296_q(16);
   n473 <= BU1296_q(15);
   n474 <= BU1296_q(14);
   n475 <= BU1296_q(13);
   n476 <= BU1296_q(12);
   n477 <= BU1296_q(11);
   n478 <= BU1296_q(10);
   n479 <= BU1296_q(9);
   n480 <= BU1296_q(8);
   n481 <= BU1296_q(7);
   n482 <= BU1296_q(6);
   n483 <= BU1296_q(5);
   n484 <= BU1296_q(4);
   n485 <= BU1296_q(3);
   n486 <= BU1296_q(2);
   n487 <= BU1296_q(1);
   n488 <= BU1296_q(0);
   BU1296_a_signed <= '0';
   BU1296_loadb <= '0';
   BU1296_swapb <= '0';
   BU1296_ce <= '1';
   BU1296_aclr <= '0';
   BU1296_sclr <= '0';
   BU1296_nd <= n341;
   n547 <= BU1296_rdy;
   BU1296 : mult_gen_v5_0
      GENERIC MAP (
         c_a_width => 14,
         c_out_width => 29,
         c_b_type => 0,
         c_has_b => 1,
         c_has_rdy => 1,
         bram_addr_width => 8,
         c_has_sclr => 0,
         c_has_nd => 1,
         c_reg_a_b_inputs => 1,
         c_enable_rlocs => 0,
         c_has_rfd => 1,
         c_mult_type => 1,
         c_has_swapb => 0,
         c_baat => 14,
         c_use_luts => 1,
         c_has_load_done => 0,
         c_has_a_signed => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 1,
         c_output_hold => 0,
         c_stack_adders => 0,
         c_mem_type => 0,
         c_b_constant => 0,
         c_has_q => 1,
         c_has_loadb => 0,
         c_pipeline => 1,
         c_has_o => 0,
         c_standalone => 1,
         c_mem_init_prefix => "mem",
         c_a_type => 0,
         c_b_width => 15,
         c_sqm_type => 0,
         c_b_value => "0"
      )
      PORT MAP (
         clk => BU1296_clk,
         a => BU1296_a,
         b => BU1296_b,
         o => BU1296_o,
         q => BU1296_q,
         a_signed => BU1296_a_signed,
         loadb => BU1296_loadb,
         load_done => BU1296_load_done,
         swapb => BU1296_swapb,
         ce => BU1296_ce,
         aclr => BU1296_aclr,
         sclr => BU1296_sclr,
         rfd => BU1296_rfd,
         nd => BU1296_nd,
         rdy => BU1296_rdy
      );

   BU1517_I(0) <= n488;
   BU1517_I(1) <= n487;
   BU1517_I(2) <= n486;
   BU1517_I(3) <= n485;
   BU1517_I(4) <= n484;
   n1547 <= BU1517_O;
   BU1517 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 5,
         c_input_inv_mask => "01111"
      )
      PORT MAP (
         I => BU1517_I,
         O => BU1517_O
      );

   BU1526_I0 <= n483;
   BU1526_I1 <= n484;
   BU1526_I2 <= n1547;
   BU1526_I3 <= '0';
   n1544 <= BU1526_O;
   BU1526 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU1526_I0,
         I1 => BU1526_I1,
         I2 => BU1526_I2,
         I3 => BU1526_I3,
         O => BU1526_O
      );

   BU1527_A(0) <= n483;
   BU1527_A(1) <= n482;
   BU1527_A(2) <= n481;
   BU1527_A(3) <= n480;
   BU1527_A(4) <= n479;
   BU1527_A(5) <= n478;
   BU1527_A(6) <= n477;
   BU1527_A(7) <= n476;
   BU1527_A(8) <= n475;
   BU1527_A(9) <= n474;
   BU1527_A(10) <= n473;
   BU1527_A(11) <= n472;
   BU1527_A(12) <= n471;
   BU1527_A(13) <= n470;
   BU1527_A(14) <= n469;
   BU1527_A(15) <= n468;
   BU1527_A(16) <= n467;
   BU1527_A(17) <= n466;
   BU1527_A(18) <= n465;
   BU1527_A(19) <= n464;
   BU1527_A(20) <= n463;
   BU1527_A(21) <= n462;
   BU1527_A(22) <= n461;
   BU1527_A(23) <= n460;
   BU1527_B(0) <= n1544;
   n1519 <= BU1527_S(0);
   n1520 <= BU1527_S(1);
   n1521 <= BU1527_S(2);
   n1522 <= BU1527_S(3);
   n1523 <= BU1527_S(4);
   n1524 <= BU1527_S(5);
   n1525 <= BU1527_S(6);
   n1526 <= BU1527_S(7);
   n1527 <= BU1527_S(8);
   n1528 <= BU1527_S(9);
   n1529 <= BU1527_S(10);
   n1530 <= BU1527_S(11);
   n1531 <= BU1527_S(12);
   n1532 <= BU1527_S(13);
   n1533 <= BU1527_S(14);
   n1534 <= BU1527_S(15);
   n1535 <= BU1527_S(16);
   n1536 <= BU1527_S(17);
   n1537 <= BU1527_S(18);
   n1538 <= BU1527_S(19);
   n1539 <= BU1527_S(20);
   n1540 <= BU1527_S(21);
   n1541 <= BU1527_S(22);
   n1542 <= BU1527_S(23);
   BU1527 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU1527_A,
         B => BU1527_B,
         S => BU1527_S
      );

   BU1628_I0 <= n460;
   BU1628_I1 <= n461;
   BU1628_I2 <= n1542;
   BU1628_I3 <= '0';
   n1553 <= BU1628_O;
   BU1628 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU1628_I0,
         I1 => BU1628_I1,
         I2 => BU1628_I2,
         I3 => BU1628_I3,
         O => BU1628_O
      );

   BU1630_I0 <= n460;
   BU1630_I1 <= n1542;
   BU1630_I2 <= '0';
   BU1630_I3 <= '0';
   n1555 <= BU1630_O;
   BU1630 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU1630_I0,
         I1 => BU1630_I1,
         I2 => BU1630_I2,
         I3 => BU1630_I3,
         O => BU1630_O
      );

   BU1631_D(0) <= n1519;
   BU1631_D(1) <= n1520;
   BU1631_D(2) <= n1521;
   BU1631_D(3) <= n1522;
   BU1631_D(4) <= n1523;
   BU1631_D(5) <= n1524;
   BU1631_D(6) <= n1525;
   BU1631_D(7) <= n1526;
   BU1631_D(8) <= n1527;
   BU1631_D(9) <= n1528;
   BU1631_D(10) <= n1529;
   BU1631_D(11) <= n1530;
   BU1631_D(12) <= n1531;
   BU1631_D(13) <= n1532;
   BU1631_D(14) <= n1533;
   BU1631_D(15) <= n1534;
   BU1631_D(16) <= n1535;
   BU1631_D(17) <= n1536;
   BU1631_D(18) <= n1537;
   BU1631_D(19) <= n1538;
   BU1631_D(20) <= n1539;
   BU1631_D(21) <= n1540;
   BU1631_D(22) <= n1541;
   n3 <= BU1631_Q(0);
   n4 <= BU1631_Q(1);
   n5 <= BU1631_Q(2);
   n6 <= BU1631_Q(3);
   n7 <= BU1631_Q(4);
   n8 <= BU1631_Q(5);
   n9 <= BU1631_Q(6);
   n10 <= BU1631_Q(7);
   n11 <= BU1631_Q(8);
   n12 <= BU1631_Q(9);
   n13 <= BU1631_Q(10);
   n14 <= BU1631_Q(11);
   n15 <= BU1631_Q(12);
   n16 <= BU1631_Q(13);
   n17 <= BU1631_Q(14);
   n18 <= BU1631_Q(15);
   n19 <= BU1631_Q(16);
   n20 <= BU1631_Q(17);
   n21 <= BU1631_Q(18);
   n22 <= BU1631_Q(19);
   n23 <= BU1631_Q(20);
   n24 <= BU1631_Q(21);
   n25 <= BU1631_Q(22);
   BU1631_CLK <= n155;
   BU1631_SCLR <= n1553;
   BU1631_SSET <= n1555;
   BU1631 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU1631_D,
         Q => BU1631_Q,
         CLK => BU1631_CLK,
         SCLR => BU1631_SCLR,
         SSET => BU1631_SSET
      );

   BU1724_D(0) <= n1542;
   n26 <= BU1724_Q(0);
   BU1724_CLK <= n155;
   BU1724_SCLR <= n1555;
   BU1724_SSET <= n1553;
   BU1724 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU1724_D,
         Q => BU1724_Q,
         CLK => BU1724_CLK,
         SCLR => BU1724_SCLR,
         SSET => BU1724_SSET
      );

   BU1729_CLK <= n155;
   BU1729_D(0) <= n547;
   n2 <= BU1729_Q(0);
   BU1729 : C_SHIFT_RAM_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_read_mif => 0,
         c_has_a => 0,
         c_sync_priority => 0,
         c_has_sclr => 0,
         c_width => 1,
         c_enable_rlocs => 0,
         c_default_data_radix => 2,
         c_generate_mif => 0,
         c_ainit_val => "0",
         c_has_ce => 0,
         c_has_aclr => 0,
         c_mem_init_radix => 2,
         c_sync_enable => 0,
         c_depth => 1,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_shift_type => 0,
         c_mem_init_file => "null",
         c_default_data => "0",
         c_reg_last_bit => 1,
         c_addr_width => 0
      )
      PORT MAP (
         CLK => BU1729_CLK,
         D => BU1729_D,
         Q => BU1729_Q
      );

   BU1734_clk <= n155;
   BU1734_a(13) <= n577;
   BU1734_a(12) <= n578;
   BU1734_a(11) <= n579;
   BU1734_a(10) <= n580;
   BU1734_a(9) <= n581;
   BU1734_a(8) <= n582;
   BU1734_a(7) <= n583;
   BU1734_a(6) <= n584;
   BU1734_a(5) <= n585;
   BU1734_a(4) <= n586;
   BU1734_a(3) <= n587;
   BU1734_a(2) <= n588;
   BU1734_a(1) <= n589;
   BU1734_a(0) <= n590;
   BU1734_b(14) <= n619;
   BU1734_b(13) <= n620;
   BU1734_b(12) <= n621;
   BU1734_b(11) <= n622;
   BU1734_b(10) <= n623;
   BU1734_b(9) <= n624;
   BU1734_b(8) <= n625;
   BU1734_b(7) <= n626;
   BU1734_b(6) <= n627;
   BU1734_b(5) <= n628;
   BU1734_b(4) <= n629;
   BU1734_b(3) <= n630;
   BU1734_b(2) <= n631;
   BU1734_b(1) <= n632;
   BU1734_b(0) <= n633;
   n664 <= BU1734_q(28);
   n665 <= BU1734_q(27);
   n666 <= BU1734_q(26);
   n667 <= BU1734_q(25);
   n668 <= BU1734_q(24);
   n669 <= BU1734_q(23);
   n670 <= BU1734_q(22);
   n671 <= BU1734_q(21);
   n672 <= BU1734_q(20);
   n673 <= BU1734_q(19);
   n674 <= BU1734_q(18);
   n675 <= BU1734_q(17);
   n676 <= BU1734_q(16);
   n677 <= BU1734_q(15);
   n678 <= BU1734_q(14);
   n679 <= BU1734_q(13);
   n680 <= BU1734_q(12);
   n681 <= BU1734_q(11);
   n682 <= BU1734_q(10);
   n683 <= BU1734_q(9);
   n684 <= BU1734_q(8);
   n685 <= BU1734_q(7);
   n686 <= BU1734_q(6);
   n687 <= BU1734_q(5);
   n688 <= BU1734_q(4);
   n689 <= BU1734_q(3);
   n690 <= BU1734_q(2);
   n691 <= BU1734_q(1);
   n692 <= BU1734_q(0);
   BU1734_a_signed <= '0';
   BU1734_loadb <= '0';
   BU1734_swapb <= '0';
   BU1734_ce <= '1';
   BU1734_aclr <= '0';
   BU1734_sclr <= '0';
   BU1734_nd <= n341;
   BU1734 : mult_gen_v5_0
      GENERIC MAP (
         c_a_width => 14,
         c_out_width => 29,
         c_b_type => 0,
         c_has_b => 1,
         c_has_rdy => 1,
         bram_addr_width => 8,
         c_has_sclr => 0,
         c_has_nd => 1,
         c_reg_a_b_inputs => 1,
         c_enable_rlocs => 0,
         c_has_rfd => 1,
         c_mult_type => 1,
         c_has_swapb => 0,
         c_baat => 14,
         c_use_luts => 1,
         c_has_load_done => 0,
         c_has_a_signed => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 1,
         c_output_hold => 0,
         c_stack_adders => 0,
         c_mem_type => 0,
         c_b_constant => 0,
         c_has_q => 1,
         c_has_loadb => 0,
         c_pipeline => 1,
         c_has_o => 0,
         c_standalone => 1,
         c_mem_init_prefix => "mem",
         c_a_type => 0,
         c_b_width => 15,
         c_sqm_type => 0,
         c_b_value => "0"
      )
      PORT MAP (
         clk => BU1734_clk,
         a => BU1734_a,
         b => BU1734_b,
         o => BU1734_o,
         q => BU1734_q,
         a_signed => BU1734_a_signed,
         loadb => BU1734_loadb,
         load_done => BU1734_load_done,
         swapb => BU1734_swapb,
         ce => BU1734_ce,
         aclr => BU1734_aclr,
         sclr => BU1734_sclr,
         rfd => BU1734_rfd,
         nd => BU1734_nd,
         rdy => BU1734_rdy
      );

   BU1955_I(0) <= n692;
   BU1955_I(1) <= n691;
   BU1955_I(2) <= n690;
   BU1955_I(3) <= n689;
   BU1955_I(4) <= n688;
   n2190 <= BU1955_O;
   BU1955 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 5,
         c_input_inv_mask => "01111"
      )
      PORT MAP (
         I => BU1955_I,
         O => BU1955_O
      );

   BU1964_I0 <= n687;
   BU1964_I1 <= n688;
   BU1964_I2 <= n2190;
   BU1964_I3 <= '0';
   n2187 <= BU1964_O;
   BU1964 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU1964_I0,
         I1 => BU1964_I1,
         I2 => BU1964_I2,
         I3 => BU1964_I3,
         O => BU1964_O
      );

   BU1965_A(0) <= n687;
   BU1965_A(1) <= n686;
   BU1965_A(2) <= n685;
   BU1965_A(3) <= n684;
   BU1965_A(4) <= n683;
   BU1965_A(5) <= n682;
   BU1965_A(6) <= n681;
   BU1965_A(7) <= n680;
   BU1965_A(8) <= n679;
   BU1965_A(9) <= n678;
   BU1965_A(10) <= n677;
   BU1965_A(11) <= n676;
   BU1965_A(12) <= n675;
   BU1965_A(13) <= n674;
   BU1965_A(14) <= n673;
   BU1965_A(15) <= n672;
   BU1965_A(16) <= n671;
   BU1965_A(17) <= n670;
   BU1965_A(18) <= n669;
   BU1965_A(19) <= n668;
   BU1965_A(20) <= n667;
   BU1965_A(21) <= n666;
   BU1965_A(22) <= n665;
   BU1965_A(23) <= n664;
   BU1965_B(0) <= n2187;
   n2162 <= BU1965_S(0);
   n2163 <= BU1965_S(1);
   n2164 <= BU1965_S(2);
   n2165 <= BU1965_S(3);
   n2166 <= BU1965_S(4);
   n2167 <= BU1965_S(5);
   n2168 <= BU1965_S(6);
   n2169 <= BU1965_S(7);
   n2170 <= BU1965_S(8);
   n2171 <= BU1965_S(9);
   n2172 <= BU1965_S(10);
   n2173 <= BU1965_S(11);
   n2174 <= BU1965_S(12);
   n2175 <= BU1965_S(13);
   n2176 <= BU1965_S(14);
   n2177 <= BU1965_S(15);
   n2178 <= BU1965_S(16);
   n2179 <= BU1965_S(17);
   n2180 <= BU1965_S(18);
   n2181 <= BU1965_S(19);
   n2182 <= BU1965_S(20);
   n2183 <= BU1965_S(21);
   n2184 <= BU1965_S(22);
   n2185 <= BU1965_S(23);
   BU1965 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU1965_A,
         B => BU1965_B,
         S => BU1965_S
      );

   BU2066_I0 <= n664;
   BU2066_I1 <= n665;
   BU2066_I2 <= n2185;
   BU2066_I3 <= '0';
   n2196 <= BU2066_O;
   BU2066 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU2066_I0,
         I1 => BU2066_I1,
         I2 => BU2066_I2,
         I3 => BU2066_I3,
         O => BU2066_O
      );

   BU2068_I0 <= n664;
   BU2068_I1 <= n2185;
   BU2068_I2 <= '0';
   BU2068_I3 <= '0';
   n2198 <= BU2068_O;
   BU2068 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU2068_I0,
         I1 => BU2068_I1,
         I2 => BU2068_I2,
         I3 => BU2068_I3,
         O => BU2068_O
      );

   BU2069_D(0) <= n2162;
   BU2069_D(1) <= n2163;
   BU2069_D(2) <= n2164;
   BU2069_D(3) <= n2165;
   BU2069_D(4) <= n2166;
   BU2069_D(5) <= n2167;
   BU2069_D(6) <= n2168;
   BU2069_D(7) <= n2169;
   BU2069_D(8) <= n2170;
   BU2069_D(9) <= n2171;
   BU2069_D(10) <= n2172;
   BU2069_D(11) <= n2173;
   BU2069_D(12) <= n2174;
   BU2069_D(13) <= n2175;
   BU2069_D(14) <= n2176;
   BU2069_D(15) <= n2177;
   BU2069_D(16) <= n2178;
   BU2069_D(17) <= n2179;
   BU2069_D(18) <= n2180;
   BU2069_D(19) <= n2181;
   BU2069_D(20) <= n2182;
   BU2069_D(21) <= n2183;
   BU2069_D(22) <= n2184;
   n27 <= BU2069_Q(0);
   n28 <= BU2069_Q(1);
   n29 <= BU2069_Q(2);
   n30 <= BU2069_Q(3);
   n31 <= BU2069_Q(4);
   n32 <= BU2069_Q(5);
   n33 <= BU2069_Q(6);
   n34 <= BU2069_Q(7);
   n35 <= BU2069_Q(8);
   n36 <= BU2069_Q(9);
   n37 <= BU2069_Q(10);
   n38 <= BU2069_Q(11);
   n39 <= BU2069_Q(12);
   n40 <= BU2069_Q(13);
   n41 <= BU2069_Q(14);
   n42 <= BU2069_Q(15);
   n43 <= BU2069_Q(16);
   n44 <= BU2069_Q(17);
   n45 <= BU2069_Q(18);
   n46 <= BU2069_Q(19);
   n47 <= BU2069_Q(20);
   n48 <= BU2069_Q(21);
   n49 <= BU2069_Q(22);
   BU2069_CLK <= n155;
   BU2069_SCLR <= n2196;
   BU2069_SSET <= n2198;
   BU2069 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2069_D,
         Q => BU2069_Q,
         CLK => BU2069_CLK,
         SCLR => BU2069_SCLR,
         SSET => BU2069_SSET
      );

   BU2162_D(0) <= n2185;
   n50 <= BU2162_Q(0);
   BU2162_CLK <= n155;
   BU2162_SCLR <= n2198;
   BU2162_SSET <= n2196;
   BU2162 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2162_D,
         Q => BU2162_Q,
         CLK => BU2162_CLK,
         SCLR => BU2162_SCLR,
         SSET => BU2162_SSET
      );

   BU2457_D <= n2726;
   BU2457_C <= n155;
   BU2457_CE <= '1';
   n2677 <= BU2457_Q;
   BU2457 : FDE
      PORT MAP (
         D => BU2457_D,
         C => BU2457_C,
         CE => BU2457_CE,
         Q => BU2457_Q
      );

   BU2461_I(0) <= n2679;
   BU2461_I(1) <= n2680;
   BU2461_I(2) <= n2681;
   BU2461_I(3) <= n2682;
   BU2461_I(4) <= n2683;
   BU2461_I(5) <= n2684;
   BU2461_I(6) <= n2685;
   BU2461_I(7) <= n2686;
   BU2461_I(8) <= n2687;
   BU2461_I(9) <= n2688;
   BU2461_I(10) <= n2689;
   BU2461_I(11) <= n2690;
   BU2461_I(12) <= n2691;
   BU2461_I(13) <= n2692;
   BU2461_I(14) <= n2693;
   BU2461_I(15) <= n2694;
   BU2461_I(16) <= n2695;
   BU2461_I(17) <= n2696;
   BU2461_I(18) <= n2697;
   BU2461_I(19) <= n2698;
   BU2461_I(20) <= n2699;
   BU2461_I(21) <= n2700;
   BU2461_I(22) <= n2701;
   n3042 <= BU2461_O;
   BU2461 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 23,
         c_input_inv_mask => "01111111111111111111111"
      )
      PORT MAP (
         I => BU2461_I,
         O => BU2461_O
      );

   BU2489_I0 <= n2702;
   BU2489_I1 <= n2701;
   BU2489_I2 <= n3042;
   BU2489_I3 <= '0';
   n3039 <= BU2489_O;
   BU2489 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU2489_I0,
         I1 => BU2489_I1,
         I2 => BU2489_I2,
         I3 => BU2489_I3,
         O => BU2489_O
      );

   BU2490_A(0) <= n2702;
   BU2490_A(1) <= n2703;
   BU2490_A(2) <= n2704;
   BU2490_A(3) <= n2705;
   BU2490_A(4) <= n2706;
   BU2490_A(5) <= n2707;
   BU2490_A(6) <= n2708;
   BU2490_A(7) <= n2709;
   BU2490_A(8) <= n2710;
   BU2490_A(9) <= n2711;
   BU2490_A(10) <= n2712;
   BU2490_A(11) <= n2713;
   BU2490_A(12) <= n2714;
   BU2490_A(13) <= n2715;
   BU2490_A(14) <= n2716;
   BU2490_A(15) <= n2717;
   BU2490_A(16) <= n2718;
   BU2490_A(17) <= n2719;
   BU2490_A(18) <= n2720;
   BU2490_A(19) <= n2721;
   BU2490_A(20) <= n2722;
   BU2490_A(21) <= n2723;
   BU2490_A(22) <= n2724;
   BU2490_A(23) <= n2725;
   BU2490_B(0) <= n3039;
   n3014 <= BU2490_S(0);
   n3015 <= BU2490_S(1);
   n3016 <= BU2490_S(2);
   n3017 <= BU2490_S(3);
   n3018 <= BU2490_S(4);
   n3019 <= BU2490_S(5);
   n3020 <= BU2490_S(6);
   n3021 <= BU2490_S(7);
   n3022 <= BU2490_S(8);
   n3023 <= BU2490_S(9);
   n3024 <= BU2490_S(10);
   n3025 <= BU2490_S(11);
   n3026 <= BU2490_S(12);
   n3027 <= BU2490_S(13);
   n3028 <= BU2490_S(14);
   n3029 <= BU2490_S(15);
   n3030 <= BU2490_S(16);
   n3031 <= BU2490_S(17);
   n3032 <= BU2490_S(18);
   n3033 <= BU2490_S(19);
   n3034 <= BU2490_S(20);
   n3035 <= BU2490_S(21);
   n3036 <= BU2490_S(22);
   n3037 <= BU2490_S(23);
   BU2490 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU2490_A,
         B => BU2490_B,
         S => BU2490_S
      );

   BU2591_I0 <= n2725;
   BU2591_I1 <= n2724;
   BU2591_I2 <= n3037;
   BU2591_I3 <= '0';
   n3066 <= BU2591_O;
   BU2591 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU2591_I0,
         I1 => BU2591_I1,
         I2 => BU2591_I2,
         I3 => BU2591_I3,
         O => BU2591_O
      );

   BU2593_I0 <= n2725;
   BU2593_I1 <= n3037;
   BU2593_I2 <= '0';
   BU2593_I3 <= '0';
   n3068 <= BU2593_O;
   BU2593 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU2593_I0,
         I1 => BU2593_I1,
         I2 => BU2593_I2,
         I3 => BU2593_I3,
         O => BU2593_O
      );

   BU2594_D(0) <= n3014;
   BU2594_D(1) <= n3015;
   BU2594_D(2) <= n3016;
   BU2594_D(3) <= n3017;
   BU2594_D(4) <= n3018;
   BU2594_D(5) <= n3019;
   BU2594_D(6) <= n3020;
   BU2594_D(7) <= n3021;
   BU2594_D(8) <= n3022;
   BU2594_D(9) <= n3023;
   BU2594_D(10) <= n3024;
   BU2594_D(11) <= n3025;
   BU2594_D(12) <= n3026;
   BU2594_D(13) <= n3027;
   BU2594_D(14) <= n3028;
   BU2594_D(15) <= n3029;
   BU2594_D(16) <= n3030;
   BU2594_D(17) <= n3031;
   BU2594_D(18) <= n3032;
   BU2594_D(19) <= n3033;
   BU2594_D(20) <= n3034;
   BU2594_D(21) <= n3035;
   BU2594_D(22) <= n3036;
   n2605 <= BU2594_Q(0);
   n2606 <= BU2594_Q(1);
   n2607 <= BU2594_Q(2);
   n2608 <= BU2594_Q(3);
   n2609 <= BU2594_Q(4);
   n2610 <= BU2594_Q(5);
   n2611 <= BU2594_Q(6);
   n2612 <= BU2594_Q(7);
   n2613 <= BU2594_Q(8);
   n2614 <= BU2594_Q(9);
   n2615 <= BU2594_Q(10);
   n2616 <= BU2594_Q(11);
   n2617 <= BU2594_Q(12);
   n2618 <= BU2594_Q(13);
   n2619 <= BU2594_Q(14);
   n2620 <= BU2594_Q(15);
   n2621 <= BU2594_Q(16);
   n2622 <= BU2594_Q(17);
   n2623 <= BU2594_Q(18);
   n2624 <= BU2594_Q(19);
   n2625 <= BU2594_Q(20);
   n2626 <= BU2594_Q(21);
   n2627 <= BU2594_Q(22);
   BU2594_CLK <= n155;
   BU2594_SCLR <= n3066;
   BU2594_SSET <= n3068;
   BU2594 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2594_D,
         Q => BU2594_Q,
         CLK => BU2594_CLK,
         SCLR => BU2594_SCLR,
         SSET => BU2594_SSET
      );

   BU2687_D(0) <= n3037;
   n2628 <= BU2687_Q(0);
   BU2687_CLK <= n155;
   BU2687_SCLR <= n3068;
   BU2687_SSET <= n3066;
   BU2687 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2687_D,
         Q => BU2687_Q,
         CLK => BU2687_CLK,
         SCLR => BU2687_SCLR,
         SSET => BU2687_SSET
      );

   BU7487_I(0) <= n2727;
   BU7487_I(1) <= n2728;
   BU7487_I(2) <= n2729;
   BU7487_I(3) <= n2730;
   BU7487_I(4) <= n2731;
   BU7487_I(5) <= n2732;
   BU7487_I(6) <= n2733;
   BU7487_I(7) <= n2734;
   BU7487_I(8) <= n2735;
   BU7487_I(9) <= n2736;
   BU7487_I(10) <= n2737;
   BU7487_I(11) <= n2738;
   BU7487_I(12) <= n2739;
   BU7487_I(13) <= n2740;
   BU7487_I(14) <= n2741;
   BU7487_I(15) <= n2742;
   BU7487_I(16) <= n2743;
   BU7487_I(17) <= n2744;
   BU7487_I(18) <= n2745;
   BU7487_I(19) <= n2746;
   BU7487_I(20) <= n2747;
   BU7487_I(21) <= n2748;
   BU7487_I(22) <= n2749;
   n3559 <= BU7487_O;
   BU7487 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 23,
         c_input_inv_mask => "01111111111111111111111"
      )
      PORT MAP (
         I => BU7487_I,
         O => BU7487_O
      );

   BU7515_I0 <= n2750;
   BU7515_I1 <= n2749;
   BU7515_I2 <= n3559;
   BU7515_I3 <= '0';
   n3556 <= BU7515_O;
   BU7515 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU7515_I0,
         I1 => BU7515_I1,
         I2 => BU7515_I2,
         I3 => BU7515_I3,
         O => BU7515_O
      );

   BU7516_A(0) <= n2750;
   BU7516_A(1) <= n2751;
   BU7516_A(2) <= n2752;
   BU7516_A(3) <= n2753;
   BU7516_A(4) <= n2754;
   BU7516_A(5) <= n2755;
   BU7516_A(6) <= n2756;
   BU7516_A(7) <= n2757;
   BU7516_A(8) <= n2758;
   BU7516_A(9) <= n2759;
   BU7516_A(10) <= n2760;
   BU7516_A(11) <= n2761;
   BU7516_A(12) <= n2762;
   BU7516_A(13) <= n2763;
   BU7516_A(14) <= n2764;
   BU7516_A(15) <= n2765;
   BU7516_A(16) <= n2766;
   BU7516_A(17) <= n2767;
   BU7516_A(18) <= n2768;
   BU7516_A(19) <= n2769;
   BU7516_A(20) <= n2770;
   BU7516_A(21) <= n2771;
   BU7516_A(22) <= n2772;
   BU7516_A(23) <= n2773;
   BU7516_B(0) <= n3556;
   n3531 <= BU7516_S(0);
   n3532 <= BU7516_S(1);
   n3533 <= BU7516_S(2);
   n3534 <= BU7516_S(3);
   n3535 <= BU7516_S(4);
   n3536 <= BU7516_S(5);
   n3537 <= BU7516_S(6);
   n3538 <= BU7516_S(7);
   n3539 <= BU7516_S(8);
   n3540 <= BU7516_S(9);
   n3541 <= BU7516_S(10);
   n3542 <= BU7516_S(11);
   n3543 <= BU7516_S(12);
   n3544 <= BU7516_S(13);
   n3545 <= BU7516_S(14);
   n3546 <= BU7516_S(15);
   n3547 <= BU7516_S(16);
   n3548 <= BU7516_S(17);
   n3549 <= BU7516_S(18);
   n3550 <= BU7516_S(19);
   n3551 <= BU7516_S(20);
   n3552 <= BU7516_S(21);
   n3553 <= BU7516_S(22);
   n3554 <= BU7516_S(23);
   BU7516 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU7516_A,
         B => BU7516_B,
         S => BU7516_S
      );

   BU7617_I0 <= n2773;
   BU7617_I1 <= n2772;
   BU7617_I2 <= n3554;
   BU7617_I3 <= '0';
   n3583 <= BU7617_O;
   BU7617 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU7617_I0,
         I1 => BU7617_I1,
         I2 => BU7617_I2,
         I3 => BU7617_I3,
         O => BU7617_O
      );

   BU7619_I0 <= n2773;
   BU7619_I1 <= n3554;
   BU7619_I2 <= '0';
   BU7619_I3 <= '0';
   n3585 <= BU7619_O;
   BU7619 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU7619_I0,
         I1 => BU7619_I1,
         I2 => BU7619_I2,
         I3 => BU7619_I3,
         O => BU7619_O
      );

   BU7620_D(0) <= n3531;
   BU7620_D(1) <= n3532;
   BU7620_D(2) <= n3533;
   BU7620_D(3) <= n3534;
   BU7620_D(4) <= n3535;
   BU7620_D(5) <= n3536;
   BU7620_D(6) <= n3537;
   BU7620_D(7) <= n3538;
   BU7620_D(8) <= n3539;
   BU7620_D(9) <= n3540;
   BU7620_D(10) <= n3541;
   BU7620_D(11) <= n3542;
   BU7620_D(12) <= n3543;
   BU7620_D(13) <= n3544;
   BU7620_D(14) <= n3545;
   BU7620_D(15) <= n3546;
   BU7620_D(16) <= n3547;
   BU7620_D(17) <= n3548;
   BU7620_D(18) <= n3549;
   BU7620_D(19) <= n3550;
   BU7620_D(20) <= n3551;
   BU7620_D(21) <= n3552;
   BU7620_D(22) <= n3553;
   n2629 <= BU7620_Q(0);
   n2630 <= BU7620_Q(1);
   n2631 <= BU7620_Q(2);
   n2632 <= BU7620_Q(3);
   n2633 <= BU7620_Q(4);
   n2634 <= BU7620_Q(5);
   n2635 <= BU7620_Q(6);
   n2636 <= BU7620_Q(7);
   n2637 <= BU7620_Q(8);
   n2638 <= BU7620_Q(9);
   n2639 <= BU7620_Q(10);
   n2640 <= BU7620_Q(11);
   n2641 <= BU7620_Q(12);
   n2642 <= BU7620_Q(13);
   n2643 <= BU7620_Q(14);
   n2644 <= BU7620_Q(15);
   n2645 <= BU7620_Q(16);
   n2646 <= BU7620_Q(17);
   n2647 <= BU7620_Q(18);
   n2648 <= BU7620_Q(19);
   n2649 <= BU7620_Q(20);
   n2650 <= BU7620_Q(21);
   n2651 <= BU7620_Q(22);
   BU7620_CLK <= n155;
   BU7620_SCLR <= n3583;
   BU7620_SSET <= n3585;
   BU7620 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU7620_D,
         Q => BU7620_Q,
         CLK => BU7620_CLK,
         SCLR => BU7620_SCLR,
         SSET => BU7620_SSET
      );

   BU7713_D(0) <= n3554;
   n2652 <= BU7713_Q(0);
   BU7713_CLK <= n155;
   BU7713_SCLR <= n3585;
   BU7713_SSET <= n3583;
   BU7713 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU7713_D,
         Q => BU7713_Q,
         CLK => BU7713_CLK,
         SCLR => BU7713_SCLR,
         SSET => BU7713_SSET
      );

   BU2173_D <= n2629;
   BU2173_C <= n155;
   BU2173_CE <= '1';
   n2653 <= BU2173_Q;
   BU2173 : FDE
      PORT MAP (
         D => BU2173_D,
         C => BU2173_C,
         CE => BU2173_CE,
         Q => BU2173_Q
      );

   BU2175_D <= n2630;
   BU2175_C <= n155;
   BU2175_CE <= '1';
   n2654 <= BU2175_Q;
   BU2175 : FDE
      PORT MAP (
         D => BU2175_D,
         C => BU2175_C,
         CE => BU2175_CE,
         Q => BU2175_Q
      );

   BU2177_D <= n2631;
   BU2177_C <= n155;
   BU2177_CE <= '1';
   n2655 <= BU2177_Q;
   BU2177 : FDE
      PORT MAP (
         D => BU2177_D,
         C => BU2177_C,
         CE => BU2177_CE,
         Q => BU2177_Q
      );

   BU2179_D <= n2632;
   BU2179_C <= n155;
   BU2179_CE <= '1';
   n2656 <= BU2179_Q;
   BU2179 : FDE
      PORT MAP (
         D => BU2179_D,
         C => BU2179_C,
         CE => BU2179_CE,
         Q => BU2179_Q
      );

   BU2181_D <= n2633;
   BU2181_C <= n155;
   BU2181_CE <= '1';
   n2657 <= BU2181_Q;
   BU2181 : FDE
      PORT MAP (
         D => BU2181_D,
         C => BU2181_C,
         CE => BU2181_CE,
         Q => BU2181_Q
      );

   BU2183_D <= n2634;
   BU2183_C <= n155;
   BU2183_CE <= '1';
   n2658 <= BU2183_Q;
   BU2183 : FDE
      PORT MAP (
         D => BU2183_D,
         C => BU2183_C,
         CE => BU2183_CE,
         Q => BU2183_Q
      );

   BU2185_D <= n2635;
   BU2185_C <= n155;
   BU2185_CE <= '1';
   n2659 <= BU2185_Q;
   BU2185 : FDE
      PORT MAP (
         D => BU2185_D,
         C => BU2185_C,
         CE => BU2185_CE,
         Q => BU2185_Q
      );

   BU2187_D <= n2636;
   BU2187_C <= n155;
   BU2187_CE <= '1';
   n2660 <= BU2187_Q;
   BU2187 : FDE
      PORT MAP (
         D => BU2187_D,
         C => BU2187_C,
         CE => BU2187_CE,
         Q => BU2187_Q
      );

   BU2189_D <= n2637;
   BU2189_C <= n155;
   BU2189_CE <= '1';
   n2661 <= BU2189_Q;
   BU2189 : FDE
      PORT MAP (
         D => BU2189_D,
         C => BU2189_C,
         CE => BU2189_CE,
         Q => BU2189_Q
      );

   BU2191_D <= n2638;
   BU2191_C <= n155;
   BU2191_CE <= '1';
   n2662 <= BU2191_Q;
   BU2191 : FDE
      PORT MAP (
         D => BU2191_D,
         C => BU2191_C,
         CE => BU2191_CE,
         Q => BU2191_Q
      );

   BU2193_D <= n2639;
   BU2193_C <= n155;
   BU2193_CE <= '1';
   n2663 <= BU2193_Q;
   BU2193 : FDE
      PORT MAP (
         D => BU2193_D,
         C => BU2193_C,
         CE => BU2193_CE,
         Q => BU2193_Q
      );

   BU2195_D <= n2640;
   BU2195_C <= n155;
   BU2195_CE <= '1';
   n2664 <= BU2195_Q;
   BU2195 : FDE
      PORT MAP (
         D => BU2195_D,
         C => BU2195_C,
         CE => BU2195_CE,
         Q => BU2195_Q
      );

   BU2197_D <= n2641;
   BU2197_C <= n155;
   BU2197_CE <= '1';
   n2665 <= BU2197_Q;
   BU2197 : FDE
      PORT MAP (
         D => BU2197_D,
         C => BU2197_C,
         CE => BU2197_CE,
         Q => BU2197_Q
      );

   BU2199_D <= n2642;
   BU2199_C <= n155;
   BU2199_CE <= '1';
   n2666 <= BU2199_Q;
   BU2199 : FDE
      PORT MAP (
         D => BU2199_D,
         C => BU2199_C,
         CE => BU2199_CE,
         Q => BU2199_Q
      );

   BU2201_D <= n2643;
   BU2201_C <= n155;
   BU2201_CE <= '1';
   n2667 <= BU2201_Q;
   BU2201 : FDE
      PORT MAP (
         D => BU2201_D,
         C => BU2201_C,
         CE => BU2201_CE,
         Q => BU2201_Q
      );

   BU2203_D <= n2644;
   BU2203_C <= n155;
   BU2203_CE <= '1';
   n2668 <= BU2203_Q;
   BU2203 : FDE
      PORT MAP (
         D => BU2203_D,
         C => BU2203_C,
         CE => BU2203_CE,
         Q => BU2203_Q
      );

   BU2205_D <= n2645;
   BU2205_C <= n155;
   BU2205_CE <= '1';
   n2669 <= BU2205_Q;
   BU2205 : FDE
      PORT MAP (
         D => BU2205_D,
         C => BU2205_C,
         CE => BU2205_CE,
         Q => BU2205_Q
      );

   BU2207_D <= n2646;
   BU2207_C <= n155;
   BU2207_CE <= '1';
   n2670 <= BU2207_Q;
   BU2207 : FDE
      PORT MAP (
         D => BU2207_D,
         C => BU2207_C,
         CE => BU2207_CE,
         Q => BU2207_Q
      );

   BU2209_D <= n2647;
   BU2209_C <= n155;
   BU2209_CE <= '1';
   n2671 <= BU2209_Q;
   BU2209 : FDE
      PORT MAP (
         D => BU2209_D,
         C => BU2209_C,
         CE => BU2209_CE,
         Q => BU2209_Q
      );

   BU2211_D <= n2648;
   BU2211_C <= n155;
   BU2211_CE <= '1';
   n2672 <= BU2211_Q;
   BU2211 : FDE
      PORT MAP (
         D => BU2211_D,
         C => BU2211_C,
         CE => BU2211_CE,
         Q => BU2211_Q
      );

   BU2213_D <= n2649;
   BU2213_C <= n155;
   BU2213_CE <= '1';
   n2673 <= BU2213_Q;
   BU2213 : FDE
      PORT MAP (
         D => BU2213_D,
         C => BU2213_C,
         CE => BU2213_CE,
         Q => BU2213_Q
      );

   BU2215_D <= n2650;
   BU2215_C <= n155;
   BU2215_CE <= '1';
   n2674 <= BU2215_Q;
   BU2215 : FDE
      PORT MAP (
         D => BU2215_D,
         C => BU2215_C,
         CE => BU2215_CE,
         Q => BU2215_Q
      );

   BU2217_D <= n2651;
   BU2217_C <= n155;
   BU2217_CE <= '1';
   n2675 <= BU2217_Q;
   BU2217 : FDE
      PORT MAP (
         D => BU2217_D,
         C => BU2217_C,
         CE => BU2217_CE,
         Q => BU2217_Q
      );

   BU2219_D <= n2652;
   BU2219_C <= n155;
   BU2219_CE <= '1';
   n2676 <= BU2219_Q;
   BU2219 : FDE
      PORT MAP (
         D => BU2219_D,
         C => BU2219_C,
         CE => BU2219_CE,
         Q => BU2219_Q
      );

   BU2220_MA(0) <= n2653;
   BU2220_MA(1) <= n2654;
   BU2220_MA(2) <= n2655;
   BU2220_MA(3) <= n2656;
   BU2220_MA(4) <= n2657;
   BU2220_MA(5) <= n2658;
   BU2220_MA(6) <= n2659;
   BU2220_MA(7) <= n2660;
   BU2220_MA(8) <= n2661;
   BU2220_MA(9) <= n2662;
   BU2220_MA(10) <= n2663;
   BU2220_MA(11) <= n2664;
   BU2220_MA(12) <= n2665;
   BU2220_MA(13) <= n2666;
   BU2220_MA(14) <= n2667;
   BU2220_MA(15) <= n2668;
   BU2220_MA(16) <= n2669;
   BU2220_MA(17) <= n2670;
   BU2220_MA(18) <= n2671;
   BU2220_MA(19) <= n2672;
   BU2220_MA(20) <= n2673;
   BU2220_MA(21) <= n2674;
   BU2220_MA(22) <= n2675;
   BU2220_MA(23) <= n2676;
   BU2220_MB(0) <= n2605;
   BU2220_MB(1) <= n2606;
   BU2220_MB(2) <= n2607;
   BU2220_MB(3) <= n2608;
   BU2220_MB(4) <= n2609;
   BU2220_MB(5) <= n2610;
   BU2220_MB(6) <= n2611;
   BU2220_MB(7) <= n2612;
   BU2220_MB(8) <= n2613;
   BU2220_MB(9) <= n2614;
   BU2220_MB(10) <= n2615;
   BU2220_MB(11) <= n2616;
   BU2220_MB(12) <= n2617;
   BU2220_MB(13) <= n2618;
   BU2220_MB(14) <= n2619;
   BU2220_MB(15) <= n2620;
   BU2220_MB(16) <= n2621;
   BU2220_MB(17) <= n2622;
   BU2220_MB(18) <= n2623;
   BU2220_MB(19) <= n2624;
   BU2220_MB(20) <= n2625;
   BU2220_MB(21) <= n2626;
   BU2220_MB(22) <= n2627;
   BU2220_MB(23) <= n2628;
   BU2220_S(0) <= n2677;
   n58 <= BU2220_Q(0);
   n59 <= BU2220_Q(1);
   n60 <= BU2220_Q(2);
   n61 <= BU2220_Q(3);
   n62 <= BU2220_Q(4);
   n63 <= BU2220_Q(5);
   n64 <= BU2220_Q(6);
   n65 <= BU2220_Q(7);
   n66 <= BU2220_Q(8);
   n67 <= BU2220_Q(9);
   n68 <= BU2220_Q(10);
   n69 <= BU2220_Q(11);
   n70 <= BU2220_Q(12);
   n71 <= BU2220_Q(13);
   n72 <= BU2220_Q(14);
   n73 <= BU2220_Q(15);
   n74 <= BU2220_Q(16);
   n75 <= BU2220_Q(17);
   n76 <= BU2220_Q(18);
   n77 <= BU2220_Q(19);
   n78 <= BU2220_Q(20);
   n79 <= BU2220_Q(21);
   n80 <= BU2220_Q(22);
   n81 <= BU2220_Q(23);
   BU2220_CLK <= n155;
   BU2220 : C_MUX_BUS_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_has_en => 0,
         c_sync_priority => 0,
         c_has_sclr => 0,
         c_width => 24,
         c_enable_rlocs => 0,
         c_sel_width => 1,
         c_latency => 1,
         c_ainit_val => "000000000000000000000000",
         c_has_ce => 0,
         c_mux_type => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "000000000000000000000000",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 1,
         c_has_o => 0,
         c_inputs => 2
      )
      PORT MAP (
         MA => BU2220_MA,
         MB => BU2220_MB,
         S => BU2220_S,
         Q => BU2220_Q,
         CLK => BU2220_CLK
      );

   BU2448_D <= n2677;
   BU2448_C <= n155;
   BU2448_CE <= '1';
   n2678 <= BU2448_Q;
   BU2448 : FDE
      PORT MAP (
         D => BU2448_D,
         C => BU2448_C,
         CE => BU2448_CE,
         Q => BU2448_Q
      );

   BU2452_I0 <= n2677;
   BU2452_I1 <= n2678;
   BU2452_I2 <= '0';
   BU2452_I3 <= '0';
   n4445 <= BU2452_O;
   BU2452 : LUT4
      GENERIC MAP (
         INIT  => X"eeee"
      )
      PORT MAP (
         I0 => BU2452_I0,
         I1 => BU2452_I1,
         I2 => BU2452_I2,
         I3 => BU2452_I3,
         O => BU2452_O
      );

   BU2453_D <= n4445;
   BU2453_C <= n155;
   BU2453_CE <= '1';
   n55 <= BU2453_Q;
   BU2453 : FDE
      PORT MAP (
         D => BU2453_D,
         C => BU2453_C,
         CE => BU2453_CE,
         Q => BU2453_Q
      );

   BU2692_DIN(0) <= n3;
   BU2692_DIN(1) <= n4;
   BU2692_DIN(2) <= n5;
   BU2692_DIN(3) <= n6;
   BU2692_DIN(4) <= n7;
   BU2692_DIN(5) <= n8;
   BU2692_DIN(6) <= n9;
   BU2692_DIN(7) <= n10;
   BU2692_DIN(8) <= n11;
   BU2692_DIN(9) <= n12;
   BU2692_DIN(10) <= n13;
   BU2692_DIN(11) <= n14;
   BU2692_DIN(12) <= n15;
   BU2692_DIN(13) <= n16;
   BU2692_DIN(14) <= n17;
   BU2692_DIN(15) <= n18;
   BU2692_DIN(16) <= n19;
   BU2692_DIN(17) <= n20;
   BU2692_DIN(18) <= n21;
   BU2692_DIN(19) <= n22;
   BU2692_DIN(20) <= n23;
   BU2692_DIN(21) <= n24;
   BU2692_DIN(22) <= n25;
   BU2692_DIN(23) <= n26;
   BU2692_ND <= n2;
   BU2692_CLK <= n155;
   n2679 <= BU2692_DOUT(0);
   n2680 <= BU2692_DOUT(1);
   n2681 <= BU2692_DOUT(2);
   n2682 <= BU2692_DOUT(3);
   n2683 <= BU2692_DOUT(4);
   n2684 <= BU2692_DOUT(5);
   n2685 <= BU2692_DOUT(6);
   n2686 <= BU2692_DOUT(7);
   n2687 <= BU2692_DOUT(8);
   n2688 <= BU2692_DOUT(9);
   n2689 <= BU2692_DOUT(10);
   n2690 <= BU2692_DOUT(11);
   n2691 <= BU2692_DOUT(12);
   n2692 <= BU2692_DOUT(13);
   n2693 <= BU2692_DOUT(14);
   n2694 <= BU2692_DOUT(15);
   n2695 <= BU2692_DOUT(16);
   n2696 <= BU2692_DOUT(17);
   n2697 <= BU2692_DOUT(18);
   n2698 <= BU2692_DOUT(19);
   n2699 <= BU2692_DOUT(20);
   n2700 <= BU2692_DOUT(21);
   n2701 <= BU2692_DOUT(22);
   n2702 <= BU2692_DOUT(23);
   n2703 <= BU2692_DOUT(24);
   n2704 <= BU2692_DOUT(25);
   n2705 <= BU2692_DOUT(26);
   n2706 <= BU2692_DOUT(27);
   n2707 <= BU2692_DOUT(28);
   n2708 <= BU2692_DOUT(29);
   n2709 <= BU2692_DOUT(30);
   n2710 <= BU2692_DOUT(31);
   n2711 <= BU2692_DOUT(32);
   n2712 <= BU2692_DOUT(33);
   n2713 <= BU2692_DOUT(34);
   n2714 <= BU2692_DOUT(35);
   n2715 <= BU2692_DOUT(36);
   n2716 <= BU2692_DOUT(37);
   n2717 <= BU2692_DOUT(38);
   n2718 <= BU2692_DOUT(39);
   n2719 <= BU2692_DOUT(40);
   n2720 <= BU2692_DOUT(41);
   n2721 <= BU2692_DOUT(42);
   n2722 <= BU2692_DOUT(43);
   n2723 <= BU2692_DOUT(44);
   n2724 <= BU2692_DOUT(45);
   n2725 <= BU2692_DOUT(46);
   n2726 <= BU2692_RDY;
   BU2692 : C_CIC_V3_0
      GENERIC MAP (
         c_differential_delay => 1,
         c_sample_rate_change_max => 16383,
         c_number_channels => 1,
         c_filter_type => 2,
         c_result_width => 47,
         c_enable_rlocs => 0,
         c_sample_rate_change => 10,
         c_latency => 1,
         c_sample_rate_change_min => 4,
         c_sample_rate_change_type => 2,
         c_data_width => 24,
         c_stages => 7
      )
      PORT MAP (
         DIN => BU2692_DIN,
         ND => BU2692_ND,
         RFD => BU2692_RFD,
         CLK => BU2692_CLK,
         DOUT => BU2692_DOUT,
         RDY => BU2692_RDY
      );

   BU7718_DIN(0) <= n27;
   BU7718_DIN(1) <= n28;
   BU7718_DIN(2) <= n29;
   BU7718_DIN(3) <= n30;
   BU7718_DIN(4) <= n31;
   BU7718_DIN(5) <= n32;
   BU7718_DIN(6) <= n33;
   BU7718_DIN(7) <= n34;
   BU7718_DIN(8) <= n35;
   BU7718_DIN(9) <= n36;
   BU7718_DIN(10) <= n37;
   BU7718_DIN(11) <= n38;
   BU7718_DIN(12) <= n39;
   BU7718_DIN(13) <= n40;
   BU7718_DIN(14) <= n41;
   BU7718_DIN(15) <= n42;
   BU7718_DIN(16) <= n43;
   BU7718_DIN(17) <= n44;
   BU7718_DIN(18) <= n45;
   BU7718_DIN(19) <= n46;
   BU7718_DIN(20) <= n47;
   BU7718_DIN(21) <= n48;
   BU7718_DIN(22) <= n49;
   BU7718_DIN(23) <= n50;
   BU7718_ND <= n2;
   BU7718_CLK <= n155;
   n2727 <= BU7718_DOUT(0);
   n2728 <= BU7718_DOUT(1);
   n2729 <= BU7718_DOUT(2);
   n2730 <= BU7718_DOUT(3);
   n2731 <= BU7718_DOUT(4);
   n2732 <= BU7718_DOUT(5);
   n2733 <= BU7718_DOUT(6);
   n2734 <= BU7718_DOUT(7);
   n2735 <= BU7718_DOUT(8);
   n2736 <= BU7718_DOUT(9);
   n2737 <= BU7718_DOUT(10);
   n2738 <= BU7718_DOUT(11);
   n2739 <= BU7718_DOUT(12);
   n2740 <= BU7718_DOUT(13);
   n2741 <= BU7718_DOUT(14);
   n2742 <= BU7718_DOUT(15);
   n2743 <= BU7718_DOUT(16);
   n2744 <= BU7718_DOUT(17);
   n2745 <= BU7718_DOUT(18);
   n2746 <= BU7718_DOUT(19);
   n2747 <= BU7718_DOUT(20);
   n2748 <= BU7718_DOUT(21);
   n2749 <= BU7718_DOUT(22);
   n2750 <= BU7718_DOUT(23);
   n2751 <= BU7718_DOUT(24);
   n2752 <= BU7718_DOUT(25);
   n2753 <= BU7718_DOUT(26);
   n2754 <= BU7718_DOUT(27);
   n2755 <= BU7718_DOUT(28);
   n2756 <= BU7718_DOUT(29);
   n2757 <= BU7718_DOUT(30);
   n2758 <= BU7718_DOUT(31);
   n2759 <= BU7718_DOUT(32);
   n2760 <= BU7718_DOUT(33);
   n2761 <= BU7718_DOUT(34);
   n2762 <= BU7718_DOUT(35);
   n2763 <= BU7718_DOUT(36);
   n2764 <= BU7718_DOUT(37);
   n2765 <= BU7718_DOUT(38);
   n2766 <= BU7718_DOUT(39);
   n2767 <= BU7718_DOUT(40);
   n2768 <= BU7718_DOUT(41);
   n2769 <= BU7718_DOUT(42);
   n2770 <= BU7718_DOUT(43);
   n2771 <= BU7718_DOUT(44);
   n2772 <= BU7718_DOUT(45);
   n2773 <= BU7718_DOUT(46);
   BU7718 : C_CIC_V3_0
      GENERIC MAP (
         c_differential_delay => 1,
         c_sample_rate_change_max => 16383,
         c_number_channels => 1,
         c_filter_type => 2,
         c_result_width => 47,
         c_enable_rlocs => 0,
         c_sample_rate_change => 10,
         c_latency => 1,
         c_sample_rate_change_min => 4,
         c_sample_rate_change_type => 2,
         c_data_width => 24,
         c_stages => 7
      )
      PORT MAP (
         DIN => BU7718_DIN,
         ND => BU7718_ND,
         RFD => BU7718_RFD,
         CLK => BU7718_CLK,
         DOUT => BU7718_DOUT,
         RDY => BU7718_RDY
      );

   BU12513_I0 <= n6719;
   BU12513_I1 <= n6691;
   BU12513_I2 <= '0';
   BU12513_I3 <= '0';
   n6718 <= BU12513_O;
   BU12513 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU12513_I0,
         I1 => BU12513_I1,
         I2 => BU12513_I2,
         I3 => BU12513_I3,
         O => BU12513_O
      );

   BU12518_I0 <= n55;
   BU12518_I1 <= '1';
   BU12518_I2 <= '0';
   BU12518_I3 <= '0';
   n6819 <= BU12518_O;
   BU12518 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU12518_I0,
         I1 => BU12518_I1,
         I2 => BU12518_I2,
         I3 => BU12518_I3,
         O => BU12518_O
      );

   BU12524_D <= '0';
   BU12524_CE <= n6819;
   BU12524_CLK <= n155;
   BU12524_A0 <= n6815;
   BU12524_A1 <= n6816;
   BU12524_A2 <= n6817;
   BU12524_A3 <= n6818;
   n6692 <= BU12524_Q;
   BU12524 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12524_D,
         CE => BU12524_CE,
         CLK => BU12524_CLK,
         A0 => BU12524_A0,
         A1 => BU12524_A1,
         A2 => BU12524_A2,
         A3 => BU12524_A3,
         Q => BU12524_Q
      );

   BU12525_D <= '0';
   BU12525_CE <= n6819;
   BU12525_CLK <= n155;
   BU12525_A0 <= n6815;
   BU12525_A1 <= n6816;
   BU12525_A2 <= n6817;
   BU12525_A3 <= n6818;
   n6693 <= BU12525_Q;
   BU12525 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12525_D,
         CE => BU12525_CE,
         CLK => BU12525_CLK,
         A0 => BU12525_A0,
         A1 => BU12525_A1,
         A2 => BU12525_A2,
         A3 => BU12525_A3,
         Q => BU12525_Q
      );

   BU12526_D <= n58;
   BU12526_CE <= n6819;
   BU12526_CLK <= n155;
   BU12526_A0 <= n6815;
   BU12526_A1 <= n6816;
   BU12526_A2 <= n6817;
   BU12526_A3 <= n6818;
   n6694 <= BU12526_Q;
   BU12526 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12526_D,
         CE => BU12526_CE,
         CLK => BU12526_CLK,
         A0 => BU12526_A0,
         A1 => BU12526_A1,
         A2 => BU12526_A2,
         A3 => BU12526_A3,
         Q => BU12526_Q
      );

   BU12527_D <= n59;
   BU12527_CE <= n6819;
   BU12527_CLK <= n155;
   BU12527_A0 <= n6815;
   BU12527_A1 <= n6816;
   BU12527_A2 <= n6817;
   BU12527_A3 <= n6818;
   n6695 <= BU12527_Q;
   BU12527 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12527_D,
         CE => BU12527_CE,
         CLK => BU12527_CLK,
         A0 => BU12527_A0,
         A1 => BU12527_A1,
         A2 => BU12527_A2,
         A3 => BU12527_A3,
         Q => BU12527_Q
      );

   BU12528_D <= n60;
   BU12528_CE <= n6819;
   BU12528_CLK <= n155;
   BU12528_A0 <= n6815;
   BU12528_A1 <= n6816;
   BU12528_A2 <= n6817;
   BU12528_A3 <= n6818;
   n6696 <= BU12528_Q;
   BU12528 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12528_D,
         CE => BU12528_CE,
         CLK => BU12528_CLK,
         A0 => BU12528_A0,
         A1 => BU12528_A1,
         A2 => BU12528_A2,
         A3 => BU12528_A3,
         Q => BU12528_Q
      );

   BU12529_D <= n61;
   BU12529_CE <= n6819;
   BU12529_CLK <= n155;
   BU12529_A0 <= n6815;
   BU12529_A1 <= n6816;
   BU12529_A2 <= n6817;
   BU12529_A3 <= n6818;
   n6697 <= BU12529_Q;
   BU12529 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12529_D,
         CE => BU12529_CE,
         CLK => BU12529_CLK,
         A0 => BU12529_A0,
         A1 => BU12529_A1,
         A2 => BU12529_A2,
         A3 => BU12529_A3,
         Q => BU12529_Q
      );

   BU12530_D <= n62;
   BU12530_CE <= n6819;
   BU12530_CLK <= n155;
   BU12530_A0 <= n6815;
   BU12530_A1 <= n6816;
   BU12530_A2 <= n6817;
   BU12530_A3 <= n6818;
   n6698 <= BU12530_Q;
   BU12530 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12530_D,
         CE => BU12530_CE,
         CLK => BU12530_CLK,
         A0 => BU12530_A0,
         A1 => BU12530_A1,
         A2 => BU12530_A2,
         A3 => BU12530_A3,
         Q => BU12530_Q
      );

   BU12531_D <= n63;
   BU12531_CE <= n6819;
   BU12531_CLK <= n155;
   BU12531_A0 <= n6815;
   BU12531_A1 <= n6816;
   BU12531_A2 <= n6817;
   BU12531_A3 <= n6818;
   n6699 <= BU12531_Q;
   BU12531 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12531_D,
         CE => BU12531_CE,
         CLK => BU12531_CLK,
         A0 => BU12531_A0,
         A1 => BU12531_A1,
         A2 => BU12531_A2,
         A3 => BU12531_A3,
         Q => BU12531_Q
      );

   BU12532_D <= n64;
   BU12532_CE <= n6819;
   BU12532_CLK <= n155;
   BU12532_A0 <= n6815;
   BU12532_A1 <= n6816;
   BU12532_A2 <= n6817;
   BU12532_A3 <= n6818;
   n6700 <= BU12532_Q;
   BU12532 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12532_D,
         CE => BU12532_CE,
         CLK => BU12532_CLK,
         A0 => BU12532_A0,
         A1 => BU12532_A1,
         A2 => BU12532_A2,
         A3 => BU12532_A3,
         Q => BU12532_Q
      );

   BU12533_D <= n65;
   BU12533_CE <= n6819;
   BU12533_CLK <= n155;
   BU12533_A0 <= n6815;
   BU12533_A1 <= n6816;
   BU12533_A2 <= n6817;
   BU12533_A3 <= n6818;
   n6701 <= BU12533_Q;
   BU12533 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12533_D,
         CE => BU12533_CE,
         CLK => BU12533_CLK,
         A0 => BU12533_A0,
         A1 => BU12533_A1,
         A2 => BU12533_A2,
         A3 => BU12533_A3,
         Q => BU12533_Q
      );

   BU12534_D <= n66;
   BU12534_CE <= n6819;
   BU12534_CLK <= n155;
   BU12534_A0 <= n6815;
   BU12534_A1 <= n6816;
   BU12534_A2 <= n6817;
   BU12534_A3 <= n6818;
   n6702 <= BU12534_Q;
   BU12534 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12534_D,
         CE => BU12534_CE,
         CLK => BU12534_CLK,
         A0 => BU12534_A0,
         A1 => BU12534_A1,
         A2 => BU12534_A2,
         A3 => BU12534_A3,
         Q => BU12534_Q
      );

   BU12535_D <= n67;
   BU12535_CE <= n6819;
   BU12535_CLK <= n155;
   BU12535_A0 <= n6815;
   BU12535_A1 <= n6816;
   BU12535_A2 <= n6817;
   BU12535_A3 <= n6818;
   n6703 <= BU12535_Q;
   BU12535 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12535_D,
         CE => BU12535_CE,
         CLK => BU12535_CLK,
         A0 => BU12535_A0,
         A1 => BU12535_A1,
         A2 => BU12535_A2,
         A3 => BU12535_A3,
         Q => BU12535_Q
      );

   BU12536_D <= n68;
   BU12536_CE <= n6819;
   BU12536_CLK <= n155;
   BU12536_A0 <= n6815;
   BU12536_A1 <= n6816;
   BU12536_A2 <= n6817;
   BU12536_A3 <= n6818;
   n6704 <= BU12536_Q;
   BU12536 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12536_D,
         CE => BU12536_CE,
         CLK => BU12536_CLK,
         A0 => BU12536_A0,
         A1 => BU12536_A1,
         A2 => BU12536_A2,
         A3 => BU12536_A3,
         Q => BU12536_Q
      );

   BU12537_D <= n69;
   BU12537_CE <= n6819;
   BU12537_CLK <= n155;
   BU12537_A0 <= n6815;
   BU12537_A1 <= n6816;
   BU12537_A2 <= n6817;
   BU12537_A3 <= n6818;
   n6705 <= BU12537_Q;
   BU12537 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12537_D,
         CE => BU12537_CE,
         CLK => BU12537_CLK,
         A0 => BU12537_A0,
         A1 => BU12537_A1,
         A2 => BU12537_A2,
         A3 => BU12537_A3,
         Q => BU12537_Q
      );

   BU12538_D <= n70;
   BU12538_CE <= n6819;
   BU12538_CLK <= n155;
   BU12538_A0 <= n6815;
   BU12538_A1 <= n6816;
   BU12538_A2 <= n6817;
   BU12538_A3 <= n6818;
   n6706 <= BU12538_Q;
   BU12538 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12538_D,
         CE => BU12538_CE,
         CLK => BU12538_CLK,
         A0 => BU12538_A0,
         A1 => BU12538_A1,
         A2 => BU12538_A2,
         A3 => BU12538_A3,
         Q => BU12538_Q
      );

   BU12539_D <= n71;
   BU12539_CE <= n6819;
   BU12539_CLK <= n155;
   BU12539_A0 <= n6815;
   BU12539_A1 <= n6816;
   BU12539_A2 <= n6817;
   BU12539_A3 <= n6818;
   n6707 <= BU12539_Q;
   BU12539 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12539_D,
         CE => BU12539_CE,
         CLK => BU12539_CLK,
         A0 => BU12539_A0,
         A1 => BU12539_A1,
         A2 => BU12539_A2,
         A3 => BU12539_A3,
         Q => BU12539_Q
      );

   BU12540_D <= n72;
   BU12540_CE <= n6819;
   BU12540_CLK <= n155;
   BU12540_A0 <= n6815;
   BU12540_A1 <= n6816;
   BU12540_A2 <= n6817;
   BU12540_A3 <= n6818;
   n6708 <= BU12540_Q;
   BU12540 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12540_D,
         CE => BU12540_CE,
         CLK => BU12540_CLK,
         A0 => BU12540_A0,
         A1 => BU12540_A1,
         A2 => BU12540_A2,
         A3 => BU12540_A3,
         Q => BU12540_Q
      );

   BU12541_D <= n73;
   BU12541_CE <= n6819;
   BU12541_CLK <= n155;
   BU12541_A0 <= n6815;
   BU12541_A1 <= n6816;
   BU12541_A2 <= n6817;
   BU12541_A3 <= n6818;
   n6709 <= BU12541_Q;
   BU12541 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12541_D,
         CE => BU12541_CE,
         CLK => BU12541_CLK,
         A0 => BU12541_A0,
         A1 => BU12541_A1,
         A2 => BU12541_A2,
         A3 => BU12541_A3,
         Q => BU12541_Q
      );

   BU12542_D <= n74;
   BU12542_CE <= n6819;
   BU12542_CLK <= n155;
   BU12542_A0 <= n6815;
   BU12542_A1 <= n6816;
   BU12542_A2 <= n6817;
   BU12542_A3 <= n6818;
   n6710 <= BU12542_Q;
   BU12542 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12542_D,
         CE => BU12542_CE,
         CLK => BU12542_CLK,
         A0 => BU12542_A0,
         A1 => BU12542_A1,
         A2 => BU12542_A2,
         A3 => BU12542_A3,
         Q => BU12542_Q
      );

   BU12543_D <= n75;
   BU12543_CE <= n6819;
   BU12543_CLK <= n155;
   BU12543_A0 <= n6815;
   BU12543_A1 <= n6816;
   BU12543_A2 <= n6817;
   BU12543_A3 <= n6818;
   n6711 <= BU12543_Q;
   BU12543 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12543_D,
         CE => BU12543_CE,
         CLK => BU12543_CLK,
         A0 => BU12543_A0,
         A1 => BU12543_A1,
         A2 => BU12543_A2,
         A3 => BU12543_A3,
         Q => BU12543_Q
      );

   BU12544_D <= n76;
   BU12544_CE <= n6819;
   BU12544_CLK <= n155;
   BU12544_A0 <= n6815;
   BU12544_A1 <= n6816;
   BU12544_A2 <= n6817;
   BU12544_A3 <= n6818;
   n6712 <= BU12544_Q;
   BU12544 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12544_D,
         CE => BU12544_CE,
         CLK => BU12544_CLK,
         A0 => BU12544_A0,
         A1 => BU12544_A1,
         A2 => BU12544_A2,
         A3 => BU12544_A3,
         Q => BU12544_Q
      );

   BU12545_D <= n77;
   BU12545_CE <= n6819;
   BU12545_CLK <= n155;
   BU12545_A0 <= n6815;
   BU12545_A1 <= n6816;
   BU12545_A2 <= n6817;
   BU12545_A3 <= n6818;
   n6713 <= BU12545_Q;
   BU12545 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12545_D,
         CE => BU12545_CE,
         CLK => BU12545_CLK,
         A0 => BU12545_A0,
         A1 => BU12545_A1,
         A2 => BU12545_A2,
         A3 => BU12545_A3,
         Q => BU12545_Q
      );

   BU12546_D <= n78;
   BU12546_CE <= n6819;
   BU12546_CLK <= n155;
   BU12546_A0 <= n6815;
   BU12546_A1 <= n6816;
   BU12546_A2 <= n6817;
   BU12546_A3 <= n6818;
   n6714 <= BU12546_Q;
   BU12546 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12546_D,
         CE => BU12546_CE,
         CLK => BU12546_CLK,
         A0 => BU12546_A0,
         A1 => BU12546_A1,
         A2 => BU12546_A2,
         A3 => BU12546_A3,
         Q => BU12546_Q
      );

   BU12547_D <= n79;
   BU12547_CE <= n6819;
   BU12547_CLK <= n155;
   BU12547_A0 <= n6815;
   BU12547_A1 <= n6816;
   BU12547_A2 <= n6817;
   BU12547_A3 <= n6818;
   n6715 <= BU12547_Q;
   BU12547 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12547_D,
         CE => BU12547_CE,
         CLK => BU12547_CLK,
         A0 => BU12547_A0,
         A1 => BU12547_A1,
         A2 => BU12547_A2,
         A3 => BU12547_A3,
         Q => BU12547_Q
      );

   BU12548_D <= n80;
   BU12548_CE <= n6819;
   BU12548_CLK <= n155;
   BU12548_A0 <= n6815;
   BU12548_A1 <= n6816;
   BU12548_A2 <= n6817;
   BU12548_A3 <= n6818;
   n6716 <= BU12548_Q;
   BU12548 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12548_D,
         CE => BU12548_CE,
         CLK => BU12548_CLK,
         A0 => BU12548_A0,
         A1 => BU12548_A1,
         A2 => BU12548_A2,
         A3 => BU12548_A3,
         Q => BU12548_Q
      );

   BU12549_D <= n81;
   BU12549_CE <= n6819;
   BU12549_CLK <= n155;
   BU12549_A0 <= n6815;
   BU12549_A1 <= n6816;
   BU12549_A2 <= n6817;
   BU12549_A3 <= n6818;
   n6717 <= BU12549_Q;
   BU12549 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12549_D,
         CE => BU12549_CE,
         CLK => BU12549_CLK,
         A0 => BU12549_A0,
         A1 => BU12549_A1,
         A2 => BU12549_A2,
         A3 => BU12549_A3,
         Q => BU12549_Q
      );

   n6815 <= BU12550_Q(0);
   n6816 <= BU12550_Q(1);
   n6817 <= BU12550_Q(2);
   n6818 <= BU12550_Q(3);
   BU12550_CLK <= n155;
   BU12550_UP <= n6819;
   BU12550_CE <= n6820;
   BU12550 : C_COUNTER_BINARY_V5_0
      GENERIC MAP (
         c_count_mode => 2,
         c_has_aset => 0,
         c_load_enable => 0,
         c_load_low => 0,
         c_count_to => "0000",
         c_sync_priority => 0,
         c_has_iv => 0,
         c_has_sclr => 0,
         c_restrict_count => 0,
         c_width => 4,
         c_has_q_thresh1 => 0,
         c_enable_rlocs => 0,
         c_has_q_thresh0 => 0,
         c_thresh1_value => "0000",
         c_has_load => 0,
         c_has_up => 0,
         c_thresh_early => 0,
         c_has_thresh1 => 0,
         c_has_thresh0 => 0,
         c_ainit_val => "0000",
         c_has_ce => 1,
         c_pipe_stages => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0000",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_count_by => "0001",
         c_has_l => 0,
         c_thresh0_value => "0000"
      )
      PORT MAP (
         Q => BU12550_Q,
         CLK => BU12550_CLK,
         UP => BU12550_UP,
         CE => BU12550_CE
      );

   BU12579_I0 <= n6718;
   BU12579_I1 <= n6819;
   BU12579_I2 <= n6719;
   BU12579_I3 <= n6821;
   n6820 <= BU12579_O;
   BU12579 : LUT4
      GENERIC MAP (
         INIT  => X"4060"
      )
      PORT MAP (
         I0 => BU12579_I0,
         I1 => BU12579_I1,
         I2 => BU12579_I2,
         I3 => BU12579_I3,
         O => BU12579_O
      );

   BU12583_I0 <= n6719;
   BU12583_I1 <= n6821;
   BU12583_I2 <= n6819;
   BU12583_I3 <= n6718;
   n7164 <= BU12583_O;
   BU12583 : LUT4
      GENERIC MAP (
         INIT  => X"e2ea"
      )
      PORT MAP (
         I0 => BU12583_I0,
         I1 => BU12583_I1,
         I2 => BU12583_I2,
         I3 => BU12583_I3,
         O => BU12583_O
      );

   BU12584_D <= n7164;
   BU12584_C <= n155;
   BU12584_CE <= '1';
   n6719 <= BU12584_Q;
   BU12584 : FDE
      PORT MAP (
         D => BU12584_D,
         C => BU12584_C,
         CE => BU12584_CE,
         Q => BU12584_Q
      );

   BU12587_I0 <= n6815;
   BU12587_I1 <= n6816;
   BU12587_I2 <= n6817;
   BU12587_I3 <= n6818;
   n6821 <= BU12587_O;
   BU12587 : LUT4
      GENERIC MAP (
         INIT  => X"0001"
      )
      PORT MAP (
         I0 => BU12587_I0,
         I1 => BU12587_I1,
         I2 => BU12587_I2,
         I3 => BU12587_I3,
         O => BU12587_O
      );

   BU12588_ND <= n6719;
   n6763 <= BU12588_RDY;
   BU12588_CLK <= n155;
   n6691 <= BU12588_RFD;
   BU12588_DIN(0) <= n6692;
   BU12588_DIN(1) <= n6693;
   BU12588_DIN(2) <= n6694;
   BU12588_DIN(3) <= n6695;
   BU12588_DIN(4) <= n6696;
   BU12588_DIN(5) <= n6697;
   BU12588_DIN(6) <= n6698;
   BU12588_DIN(7) <= n6699;
   BU12588_DIN(8) <= n6700;
   BU12588_DIN(9) <= n6701;
   BU12588_DIN(10) <= n6702;
   BU12588_DIN(11) <= n6703;
   BU12588_DIN(12) <= n6704;
   BU12588_DIN(13) <= n6705;
   BU12588_DIN(14) <= n6706;
   BU12588_DIN(15) <= n6707;
   BU12588_DIN(16) <= n6708;
   BU12588_DIN(17) <= n6709;
   BU12588_DIN(18) <= n6710;
   BU12588_DIN(19) <= n6711;
   BU12588_DIN(20) <= n6712;
   BU12588_DIN(21) <= n6713;
   BU12588_DIN(22) <= n6714;
   BU12588_DIN(23) <= n6715;
   BU12588_DIN(24) <= n6716;
   BU12588_DIN(25) <= n6717;
   n6720 <= BU12588_DOUT(0);
   n6721 <= BU12588_DOUT(1);
   n6722 <= BU12588_DOUT(2);
   n6723 <= BU12588_DOUT(3);
   n6724 <= BU12588_DOUT(4);
   n6725 <= BU12588_DOUT(5);
   n6726 <= BU12588_DOUT(6);
   n6727 <= BU12588_DOUT(7);
   n6728 <= BU12588_DOUT(8);
   n6729 <= BU12588_DOUT(9);
   n6730 <= BU12588_DOUT(10);
   n6731 <= BU12588_DOUT(11);
   n6732 <= BU12588_DOUT(12);
   n6733 <= BU12588_DOUT(13);
   n6734 <= BU12588_DOUT(14);
   n6735 <= BU12588_DOUT(15);
   n6736 <= BU12588_DOUT(16);
   n6737 <= BU12588_DOUT(17);
   n6738 <= BU12588_DOUT(18);
   n6739 <= BU12588_DOUT(19);
   n6740 <= BU12588_DOUT(20);
   n6741 <= BU12588_DOUT(21);
   n6742 <= BU12588_DOUT(22);
   n6743 <= BU12588_DOUT(23);
   n6744 <= BU12588_DOUT(24);
   n6745 <= BU12588_DOUT(25);
   n6746 <= BU12588_DOUT(26);
   n6747 <= BU12588_DOUT(27);
   n6748 <= BU12588_DOUT(28);
   n6749 <= BU12588_DOUT(29);
   n6750 <= BU12588_DOUT(30);
   n6751 <= BU12588_DOUT(31);
   n6752 <= BU12588_DOUT(32);
   n6753 <= BU12588_DOUT(33);
   n6754 <= BU12588_DOUT(34);
   n6755 <= BU12588_DOUT(35);
   n6756 <= BU12588_DOUT(36);
   n6757 <= BU12588_DOUT(37);
   n6758 <= BU12588_DOUT(38);
   n6759 <= BU12588_DOUT(39);
   n6760 <= BU12588_DOUT(40);
   n6761 <= BU12588_DOUT(41);
   n6762 <= BU12588_DOUT(42);
   BU12588 : C_DA_FIR_V7_0
      GENERIC MAP (
         c_has_sout_r => 0,
         c_result_width => 43,
         c_reload_delay => 401,
         c_data_type => 0,
         c_filter_type => 0,
         c_channels => 2,
         c_response => 0,
         c_has_sout_f => 0,
         c_reg_output => 0,
         c_taps => 45,
         c_data_width => 26,
         c_enable_rlocs => 0,
         c_coeff_type => 0,
         c_reload_mem_type => 2,
         c_has_sin_r => 0,
         c_reload => 0,
         c_baat => 6,
         c_latency => 15,
         c_coeff_width => 16,
         c_optimize => 1,
         c_use_model_func => 0,
         c_zpf => 1,
         c_has_sin_f => 0,
         c_shape => 0,
         c_saturate => 0,
         c_has_sel_o => 0,
         c_mem_init_file => "ddcv_orig_CFIR.mif",
         c_polyphase_factor => 1,
         c_has_sel_i => 0,
         c_has_reset => 0
      )
      PORT MAP (
         ND => BU12588_ND,
         RDY => BU12588_RDY,
         CLK => BU12588_CLK,
         RFD => BU12588_RFD,
         DIN => BU12588_DIN,
         DOUT => BU12588_DOUT
      );

   BU19118_I(0) <= n6720;
   BU19118_I(1) <= n6721;
   BU19118_I(2) <= n6722;
   BU19118_I(3) <= n6723;
   BU19118_I(4) <= n6724;
   BU19118_I(5) <= n6725;
   BU19118_I(6) <= n6726;
   BU19118_I(7) <= n6727;
   BU19118_I(8) <= n6728;
   BU19118_I(9) <= n6729;
   BU19118_I(10) <= n6730;
   BU19118_I(11) <= n6731;
   BU19118_I(12) <= n6732;
   BU19118_I(13) <= n6733;
   BU19118_I(14) <= n6734;
   BU19118_I(15) <= n6735;
   BU19118_I(16) <= n6736;
   BU19118_I(17) <= n6737;
   BU19118_I(18) <= n6738;
   BU19118_I(19) <= n6739;
   BU19118_I(20) <= n6740;
   BU19118_I(21) <= n6741;
   BU19118_I(22) <= n6742;
   BU19118_I(23) <= n6743;
   BU19118_I(24) <= n6744;
   BU19118_I(25) <= n6745;
   BU19118_I(26) <= n6746;
   n7297 <= BU19118_O;
   BU19118 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 27,
         c_input_inv_mask => "011111111111111111111111111"
      )
      PORT MAP (
         I => BU19118_I,
         O => BU19118_O
      );

   BU19149_I0 <= n6747;
   BU19149_I1 <= n6746;
   BU19149_I2 <= n7297;
   BU19149_I3 <= '0';
   n7294 <= BU19149_O;
   BU19149 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU19149_I0,
         I1 => BU19149_I1,
         I2 => BU19149_I2,
         I3 => BU19149_I3,
         O => BU19149_O
      );

   BU19150_A(0) <= n6747;
   BU19150_A(1) <= n6748;
   BU19150_A(2) <= n6749;
   BU19150_A(3) <= n6750;
   BU19150_A(4) <= n6751;
   BU19150_A(5) <= n6752;
   BU19150_A(6) <= n6753;
   BU19150_A(7) <= n6754;
   BU19150_A(8) <= n6755;
   BU19150_A(9) <= n6756;
   BU19150_A(10) <= n6757;
   BU19150_A(11) <= n6758;
   BU19150_A(12) <= n6759;
   BU19150_A(13) <= n6760;
   BU19150_A(14) <= n6761;
   BU19150_A(15) <= n6762;
   BU19150_B(0) <= n7294;
   n7277 <= BU19150_S(0);
   n7278 <= BU19150_S(1);
   n7279 <= BU19150_S(2);
   n7280 <= BU19150_S(3);
   n7281 <= BU19150_S(4);
   n7282 <= BU19150_S(5);
   n7283 <= BU19150_S(6);
   n7284 <= BU19150_S(7);
   n7285 <= BU19150_S(8);
   n7286 <= BU19150_S(9);
   n7287 <= BU19150_S(10);
   n7288 <= BU19150_S(11);
   n7289 <= BU19150_S(12);
   n7290 <= BU19150_S(13);
   n7291 <= BU19150_S(14);
   n7292 <= BU19150_S(15);
   BU19150 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 16,
         c_latency => 1,
         c_sinit_val => "00000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "00000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 17,
         c_low_bit => 0,
         c_ainit_val => "00000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 16,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU19150_A,
         B => BU19150_B,
         S => BU19150_S
      );

   BU19219_I0 <= n6762;
   BU19219_I1 <= n6761;
   BU19219_I2 <= n7292;
   BU19219_I3 <= '0';
   n7325 <= BU19219_O;
   BU19219 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU19219_I0,
         I1 => BU19219_I1,
         I2 => BU19219_I2,
         I3 => BU19219_I3,
         O => BU19219_O
      );

   BU19221_I0 <= n6762;
   BU19221_I1 <= n7292;
   BU19221_I2 <= '0';
   BU19221_I3 <= '0';
   n7327 <= BU19221_O;
   BU19221 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU19221_I0,
         I1 => BU19221_I1,
         I2 => BU19221_I2,
         I3 => BU19221_I3,
         O => BU19221_O
      );

   BU19222_D(0) <= n7277;
   BU19222_D(1) <= n7278;
   BU19222_D(2) <= n7279;
   BU19222_D(3) <= n7280;
   BU19222_D(4) <= n7281;
   BU19222_D(5) <= n7282;
   BU19222_D(6) <= n7283;
   BU19222_D(7) <= n7284;
   BU19222_D(8) <= n7285;
   BU19222_D(9) <= n7286;
   BU19222_D(10) <= n7287;
   BU19222_D(11) <= n7288;
   BU19222_D(12) <= n7289;
   BU19222_D(13) <= n7290;
   BU19222_D(14) <= n7291;
   n82 <= BU19222_Q(0);
   n83 <= BU19222_Q(1);
   n84 <= BU19222_Q(2);
   n85 <= BU19222_Q(3);
   n86 <= BU19222_Q(4);
   n87 <= BU19222_Q(5);
   n88 <= BU19222_Q(6);
   n89 <= BU19222_Q(7);
   n90 <= BU19222_Q(8);
   n91 <= BU19222_Q(9);
   n92 <= BU19222_Q(10);
   n93 <= BU19222_Q(11);
   n94 <= BU19222_Q(12);
   n95 <= BU19222_Q(13);
   n96 <= BU19222_Q(14);
   BU19222_CLK <= n155;
   BU19222_SCLR <= n7325;
   BU19222_SSET <= n7327;
   BU19222 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 15,
         c_has_ce => 0,
         c_sinit_val => "000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU19222_D,
         Q => BU19222_Q,
         CLK => BU19222_CLK,
         SCLR => BU19222_SCLR,
         SSET => BU19222_SSET
      );

   BU19283_D(0) <= n7292;
   n97 <= BU19283_Q(0);
   BU19283_CLK <= n155;
   BU19283_SCLR <= n7327;
   BU19283_SSET <= n7325;
   BU19283 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU19283_D,
         Q => BU19283_Q,
         CLK => BU19283_CLK,
         SCLR => BU19283_SCLR,
         SSET => BU19283_SSET
      );

   BU19290_D <= n6763;
   BU19290_C <= n155;
   BU19290_CE <= '1';
   n98 <= BU19290_Q;
   BU19290 : FDE
      PORT MAP (
         D => BU19290_D,
         C => BU19290_C,
         CE => BU19290_CE,
         Q => BU19290_Q
      );

   BU19293_ND <= n98;
   n134 <= BU19293_RDY;
   BU19293_CLK <= n155;
   BU19293_DIN(0) <= n82;
   BU19293_DIN(1) <= n83;
   BU19293_DIN(2) <= n84;
   BU19293_DIN(3) <= n85;
   BU19293_DIN(4) <= n86;
   BU19293_DIN(5) <= n87;
   BU19293_DIN(6) <= n88;
   BU19293_DIN(7) <= n89;
   BU19293_DIN(8) <= n90;
   BU19293_DIN(9) <= n91;
   BU19293_DIN(10) <= n92;
   BU19293_DIN(11) <= n93;
   BU19293_DIN(12) <= n94;
   BU19293_DIN(13) <= n95;
   BU19293_DIN(14) <= n96;
   BU19293_DIN(15) <= n97;
   n135 <= BU19293_SEL_O(0);
   n99 <= BU19293_DOUT(0);
   n100 <= BU19293_DOUT(1);
   n101 <= BU19293_DOUT(2);
   n102 <= BU19293_DOUT(3);
   n103 <= BU19293_DOUT(4);
   n104 <= BU19293_DOUT(5);
   n105 <= BU19293_DOUT(6);
   n106 <= BU19293_DOUT(7);
   n107 <= BU19293_DOUT(8);
   n108 <= BU19293_DOUT(9);
   n109 <= BU19293_DOUT(10);
   n110 <= BU19293_DOUT(11);
   n111 <= BU19293_DOUT(12);
   n112 <= BU19293_DOUT(13);
   n113 <= BU19293_DOUT(14);
   n114 <= BU19293_DOUT(15);
   n115 <= BU19293_DOUT(16);
   n116 <= BU19293_DOUT(17);
   n117 <= BU19293_DOUT(18);
   n118 <= BU19293_DOUT(19);
   n119 <= BU19293_DOUT(20);
   n120 <= BU19293_DOUT(21);
   n121 <= BU19293_DOUT(22);
   n122 <= BU19293_DOUT(23);
   n123 <= BU19293_DOUT(24);
   n124 <= BU19293_DOUT(25);
   n125 <= BU19293_DOUT(26);
   n126 <= BU19293_DOUT(27);
   n127 <= BU19293_DOUT(28);
   n128 <= BU19293_DOUT(29);
   n129 <= BU19293_DOUT(30);
   n130 <= BU19293_DOUT(31);
   n131 <= BU19293_DOUT(32);
   n132 <= BU19293_DOUT(33);
   n133 <= BU19293_DOUT(34);
   BU19293 : C_DA_FIR_V7_0
      GENERIC MAP (
         c_has_sout_r => 0,
         c_result_width => 35,
         c_reload_delay => 657,
         c_data_type => 0,
         c_filter_type => 2,
         c_channels => 2,
         c_response => 0,
         c_has_sout_f => 0,
         c_reg_output => 0,
         c_taps => 55,
         c_data_width => 16,
         c_enable_rlocs => 0,
         c_coeff_type => 0,
         c_reload_mem_type => 2,
         c_has_sin_r => 0,
         c_reload => 0,
         c_baat => 1,
         c_latency => 26,
         c_coeff_width => 16,
         c_optimize => 1,
         c_use_model_func => 0,
         c_zpf => 1,
         c_has_sin_f => 0,
         c_shape => 0,
         c_saturate => 0,
         c_has_sel_o => 1,
         c_mem_init_file => "ddcv_orig_PFIR.mif",
         c_polyphase_factor => 5,
         c_has_sel_i => 0,
         c_has_reset => 0
      )
      PORT MAP (
         ND => BU19293_ND,
         RDY => BU19293_RDY,
         CLK => BU19293_CLK,
         RFD => BU19293_RFD,
         DIN => BU19293_DIN,
         SEL_O => BU19293_SEL_O,
         DOUT => BU19293_DOUT
      );

   BU22774_I0 <= n134;
   BU22774_I1 <= n135;
   BU22774_I2 <= '0';
   BU22774_I3 <= '0';
   n136 <= BU22774_O;
   BU22774 : LUT4
      GENERIC MAP (
         INIT  => X"2222"
      )
      PORT MAP (
         I0 => BU22774_I0,
         I1 => BU22774_I1,
         I2 => BU22774_I2,
         I3 => BU22774_I3,
         O => BU22774_O
      );

   BU22776_I0 <= n134;
   BU22776_I1 <= n135;
   BU22776_I2 <= '0';
   BU22776_I3 <= '0';
   n137 <= BU22776_O;
   BU22776 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU22776_I0,
         I1 => BU22776_I1,
         I2 => BU22776_I2,
         I3 => BU22776_I3,
         O => BU22776_O
      );

   BU22779_D <= n137;
   BU22779_C <= n155;
   BU22779_CE <= '1';
   n153 <= BU22779_Q;
   BU22779 : FDE
      PORT MAP (
         D => BU22779_D,
         C => BU22779_C,
         CE => BU22779_CE,
         Q => BU22779_Q
      );

   BU22784_I(0) <= n99;
   BU22784_I(1) <= n100;
   BU22784_I(2) <= n101;
   BU22784_I(3) <= n102;
   BU22784_I(4) <= n103;
   n7868 <= BU22784_O;
   BU22784 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 5,
         c_input_inv_mask => "01111"
      )
      PORT MAP (
         I => BU22784_I,
         O => BU22784_O
      );

   BU22793_I0 <= n104;
   BU22793_I1 <= n103;
   BU22793_I2 <= n7868;
   BU22793_I3 <= '0';
   n7865 <= BU22793_O;
   BU22793 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU22793_I0,
         I1 => BU22793_I1,
         I2 => BU22793_I2,
         I3 => BU22793_I3,
         O => BU22793_O
      );

   BU22794_A(0) <= n104;
   BU22794_A(1) <= n105;
   BU22794_A(2) <= n106;
   BU22794_A(3) <= n107;
   BU22794_A(4) <= n108;
   BU22794_A(5) <= n109;
   BU22794_A(6) <= n110;
   BU22794_A(7) <= n111;
   BU22794_A(8) <= n112;
   BU22794_A(9) <= n113;
   BU22794_A(10) <= n114;
   BU22794_A(11) <= n115;
   BU22794_A(12) <= n116;
   BU22794_A(13) <= n117;
   BU22794_A(14) <= n118;
   BU22794_A(15) <= n119;
   BU22794_A(16) <= n120;
   BU22794_A(17) <= n121;
   BU22794_A(18) <= n122;
   BU22794_A(19) <= n123;
   BU22794_A(20) <= n124;
   BU22794_A(21) <= n125;
   BU22794_A(22) <= n126;
   BU22794_A(23) <= n127;
   BU22794_A(24) <= n128;
   BU22794_A(25) <= n129;
   BU22794_A(26) <= n130;
   BU22794_A(27) <= n131;
   BU22794_A(28) <= n132;
   BU22794_A(29) <= n133;
   BU22794_B(0) <= n7865;
   n7834 <= BU22794_S(0);
   n7835 <= BU22794_S(1);
   n7836 <= BU22794_S(2);
   n7837 <= BU22794_S(3);
   n7838 <= BU22794_S(4);
   n7839 <= BU22794_S(5);
   n7840 <= BU22794_S(6);
   n7841 <= BU22794_S(7);
   n7842 <= BU22794_S(8);
   n7843 <= BU22794_S(9);
   n7844 <= BU22794_S(10);
   n7845 <= BU22794_S(11);
   n7846 <= BU22794_S(12);
   n7847 <= BU22794_S(13);
   n7848 <= BU22794_S(14);
   n7849 <= BU22794_S(15);
   n7850 <= BU22794_S(16);
   n7851 <= BU22794_S(17);
   n7852 <= BU22794_S(18);
   n7853 <= BU22794_S(19);
   n7854 <= BU22794_S(20);
   n7855 <= BU22794_S(21);
   n7856 <= BU22794_S(22);
   n7857 <= BU22794_S(23);
   n7858 <= BU22794_S(24);
   n7859 <= BU22794_S(25);
   n7860 <= BU22794_S(26);
   n7861 <= BU22794_S(27);
   n7862 <= BU22794_S(28);
   n7863 <= BU22794_S(29);
   BU22794 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 30,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 31,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 30,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU22794_A,
         B => BU22794_B,
         S => BU22794_S
      );

   BU22919_I0 <= n133;
   BU22919_I1 <= n132;
   BU22919_I2 <= n7863;
   BU22919_I3 <= n136;
   n7874 <= BU22919_O;
   BU22919 : LUT4
      GENERIC MAP (
         INIT  => X"0200"
      )
      PORT MAP (
         I0 => BU22919_I0,
         I1 => BU22919_I1,
         I2 => BU22919_I2,
         I3 => BU22919_I3,
         O => BU22919_O
      );

   BU22921_I0 <= n133;
   BU22921_I1 <= n7863;
   BU22921_I2 <= n136;
   BU22921_I3 <= '0';
   n7876 <= BU22921_O;
   BU22921 : LUT4
      GENERIC MAP (
         INIT  => X"4040"
      )
      PORT MAP (
         I0 => BU22921_I0,
         I1 => BU22921_I1,
         I2 => BU22921_I2,
         I3 => BU22921_I3,
         O => BU22921_O
      );

   BU22922_D(0) <= n7834;
   BU22922_D(1) <= n7835;
   BU22922_D(2) <= n7836;
   BU22922_D(3) <= n7837;
   BU22922_D(4) <= n7838;
   BU22922_D(5) <= n7839;
   BU22922_D(6) <= n7840;
   BU22922_D(7) <= n7841;
   BU22922_D(8) <= n7842;
   BU22922_D(9) <= n7843;
   BU22922_D(10) <= n7844;
   BU22922_D(11) <= n7845;
   BU22922_D(12) <= n7846;
   BU22922_D(13) <= n7847;
   BU22922_D(14) <= n7848;
   BU22922_D(15) <= n7849;
   BU22922_D(16) <= n7850;
   BU22922_D(17) <= n7851;
   BU22922_D(18) <= n7852;
   BU22922_D(19) <= n7853;
   BU22922_D(20) <= n7854;
   BU22922_D(21) <= n7855;
   BU22922_D(22) <= n7856;
   BU22922_D(23) <= n7857;
   BU22922_D(24) <= n7858;
   BU22922_D(25) <= n7859;
   BU22922_D(26) <= n7860;
   BU22922_D(27) <= n7861;
   BU22922_D(28) <= n7862;
   n195 <= BU22922_Q(0);
   n196 <= BU22922_Q(1);
   n197 <= BU22922_Q(2);
   n198 <= BU22922_Q(3);
   n199 <= BU22922_Q(4);
   n200 <= BU22922_Q(5);
   n201 <= BU22922_Q(6);
   n202 <= BU22922_Q(7);
   n203 <= BU22922_Q(8);
   n204 <= BU22922_Q(9);
   n205 <= BU22922_Q(10);
   n206 <= BU22922_Q(11);
   n207 <= BU22922_Q(12);
   n208 <= BU22922_Q(13);
   n209 <= BU22922_Q(14);
   n210 <= BU22922_Q(15);
   n211 <= BU22922_Q(16);
   n212 <= BU22922_Q(17);
   n213 <= BU22922_Q(18);
   n214 <= BU22922_Q(19);
   n215 <= BU22922_Q(20);
   n216 <= BU22922_Q(21);
   n217 <= BU22922_Q(22);
   n218 <= BU22922_Q(23);
   n219 <= BU22922_Q(24);
   n220 <= BU22922_Q(25);
   n221 <= BU22922_Q(26);
   n222 <= BU22922_Q(27);
   n223 <= BU22922_Q(28);
   BU22922_CLK <= n155;
   BU22922_CE <= n136;
   BU22922_SCLR <= n7874;
   BU22922_SSET <= n7876;
   BU22922 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 29,
         c_has_ce => 1,
         c_sinit_val => "00000000000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU22922_D,
         Q => BU22922_Q,
         CLK => BU22922_CLK,
         CE => BU22922_CE,
         SCLR => BU22922_SCLR,
         SSET => BU22922_SSET
      );

   BU23042_D(0) <= n7863;
   n224 <= BU23042_Q(0);
   BU23042_CLK <= n155;
   BU23042_CE <= n136;
   BU23042_SCLR <= n7876;
   BU23042_SSET <= n7874;
   BU23042 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 1,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU23042_D,
         Q => BU23042_Q,
         CLK => BU23042_CLK,
         CE => BU23042_CE,
         SCLR => BU23042_SCLR,
         SSET => BU23042_SSET
      );

   BU23054_I(0) <= n99;
   BU23054_I(1) <= n100;
   BU23054_I(2) <= n101;
   BU23054_I(3) <= n102;
   BU23054_I(4) <= n103;
   n8413 <= BU23054_O;
   BU23054 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 5,
         c_input_inv_mask => "01111"
      )
      PORT MAP (
         I => BU23054_I,
         O => BU23054_O
      );

   BU23063_I0 <= n104;
   BU23063_I1 <= n103;
   BU23063_I2 <= n8413;
   BU23063_I3 <= '0';
   n8410 <= BU23063_O;
   BU23063 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU23063_I0,
         I1 => BU23063_I1,
         I2 => BU23063_I2,
         I3 => BU23063_I3,
         O => BU23063_O
      );

   BU23064_A(0) <= n104;
   BU23064_A(1) <= n105;
   BU23064_A(2) <= n106;
   BU23064_A(3) <= n107;
   BU23064_A(4) <= n108;
   BU23064_A(5) <= n109;
   BU23064_A(6) <= n110;
   BU23064_A(7) <= n111;
   BU23064_A(8) <= n112;
   BU23064_A(9) <= n113;
   BU23064_A(10) <= n114;
   BU23064_A(11) <= n115;
   BU23064_A(12) <= n116;
   BU23064_A(13) <= n117;
   BU23064_A(14) <= n118;
   BU23064_A(15) <= n119;
   BU23064_A(16) <= n120;
   BU23064_A(17) <= n121;
   BU23064_A(18) <= n122;
   BU23064_A(19) <= n123;
   BU23064_A(20) <= n124;
   BU23064_A(21) <= n125;
   BU23064_A(22) <= n126;
   BU23064_A(23) <= n127;
   BU23064_A(24) <= n128;
   BU23064_A(25) <= n129;
   BU23064_A(26) <= n130;
   BU23064_A(27) <= n131;
   BU23064_A(28) <= n132;
   BU23064_A(29) <= n133;
   BU23064_B(0) <= n8410;
   n8379 <= BU23064_S(0);
   n8380 <= BU23064_S(1);
   n8381 <= BU23064_S(2);
   n8382 <= BU23064_S(3);
   n8383 <= BU23064_S(4);
   n8384 <= BU23064_S(5);
   n8385 <= BU23064_S(6);
   n8386 <= BU23064_S(7);
   n8387 <= BU23064_S(8);
   n8388 <= BU23064_S(9);
   n8389 <= BU23064_S(10);
   n8390 <= BU23064_S(11);
   n8391 <= BU23064_S(12);
   n8392 <= BU23064_S(13);
   n8393 <= BU23064_S(14);
   n8394 <= BU23064_S(15);
   n8395 <= BU23064_S(16);
   n8396 <= BU23064_S(17);
   n8397 <= BU23064_S(18);
   n8398 <= BU23064_S(19);
   n8399 <= BU23064_S(20);
   n8400 <= BU23064_S(21);
   n8401 <= BU23064_S(22);
   n8402 <= BU23064_S(23);
   n8403 <= BU23064_S(24);
   n8404 <= BU23064_S(25);
   n8405 <= BU23064_S(26);
   n8406 <= BU23064_S(27);
   n8407 <= BU23064_S(28);
   n8408 <= BU23064_S(29);
   BU23064 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 30,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 31,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 30,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU23064_A,
         B => BU23064_B,
         S => BU23064_S
      );

   BU23189_I0 <= n133;
   BU23189_I1 <= n132;
   BU23189_I2 <= n8408;
   BU23189_I3 <= n137;
   n8419 <= BU23189_O;
   BU23189 : LUT4
      GENERIC MAP (
         INIT  => X"0200"
      )
      PORT MAP (
         I0 => BU23189_I0,
         I1 => BU23189_I1,
         I2 => BU23189_I2,
         I3 => BU23189_I3,
         O => BU23189_O
      );

   BU23191_I0 <= n133;
   BU23191_I1 <= n8408;
   BU23191_I2 <= n137;
   BU23191_I3 <= '0';
   n8421 <= BU23191_O;
   BU23191 : LUT4
      GENERIC MAP (
         INIT  => X"4040"
      )
      PORT MAP (
         I0 => BU23191_I0,
         I1 => BU23191_I1,
         I2 => BU23191_I2,
         I3 => BU23191_I3,
         O => BU23191_O
      );

   BU23192_D(0) <= n8379;
   BU23192_D(1) <= n8380;
   BU23192_D(2) <= n8381;
   BU23192_D(3) <= n8382;
   BU23192_D(4) <= n8383;
   BU23192_D(5) <= n8384;
   BU23192_D(6) <= n8385;
   BU23192_D(7) <= n8386;
   BU23192_D(8) <= n8387;
   BU23192_D(9) <= n8388;
   BU23192_D(10) <= n8389;
   BU23192_D(11) <= n8390;
   BU23192_D(12) <= n8391;
   BU23192_D(13) <= n8392;
   BU23192_D(14) <= n8393;
   BU23192_D(15) <= n8394;
   BU23192_D(16) <= n8395;
   BU23192_D(17) <= n8396;
   BU23192_D(18) <= n8397;
   BU23192_D(19) <= n8398;
   BU23192_D(20) <= n8399;
   BU23192_D(21) <= n8400;
   BU23192_D(22) <= n8401;
   BU23192_D(23) <= n8402;
   BU23192_D(24) <= n8403;
   BU23192_D(25) <= n8404;
   BU23192_D(26) <= n8405;
   BU23192_D(27) <= n8406;
   BU23192_D(28) <= n8407;
   n225 <= BU23192_Q(0);
   n226 <= BU23192_Q(1);
   n227 <= BU23192_Q(2);
   n228 <= BU23192_Q(3);
   n229 <= BU23192_Q(4);
   n230 <= BU23192_Q(5);
   n231 <= BU23192_Q(6);
   n232 <= BU23192_Q(7);
   n233 <= BU23192_Q(8);
   n234 <= BU23192_Q(9);
   n235 <= BU23192_Q(10);
   n236 <= BU23192_Q(11);
   n237 <= BU23192_Q(12);
   n238 <= BU23192_Q(13);
   n239 <= BU23192_Q(14);
   n240 <= BU23192_Q(15);
   n241 <= BU23192_Q(16);
   n242 <= BU23192_Q(17);
   n243 <= BU23192_Q(18);
   n244 <= BU23192_Q(19);
   n245 <= BU23192_Q(20);
   n246 <= BU23192_Q(21);
   n247 <= BU23192_Q(22);
   n248 <= BU23192_Q(23);
   n249 <= BU23192_Q(24);
   n250 <= BU23192_Q(25);
   n251 <= BU23192_Q(26);
   n252 <= BU23192_Q(27);
   n253 <= BU23192_Q(28);
   BU23192_CLK <= n155;
   BU23192_CE <= n137;
   BU23192_SCLR <= n8419;
   BU23192_SSET <= n8421;
   BU23192 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 29,
         c_has_ce => 1,
         c_sinit_val => "00000000000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU23192_D,
         Q => BU23192_Q,
         CLK => BU23192_CLK,
         CE => BU23192_CE,
         SCLR => BU23192_SCLR,
         SSET => BU23192_SSET
      );

   BU23312_D(0) <= n8408;
   n254 <= BU23312_Q(0);
   BU23312_CLK <= n155;
   BU23312_CE <= n137;
   BU23312_SCLR <= n8421;
   BU23312_SSET <= n8419;
   BU23312 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 1,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU23312_D,
         Q => BU23312_Q,
         CLK => BU23312_CLK,
         CE => BU23312_CE,
         SCLR => BU23312_SCLR,
         SSET => BU23312_SSET
      );


END xilinx;


-- synopsys translate_on
