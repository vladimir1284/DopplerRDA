--------------------------------------------------------------------------------
--     This file is owned and controlled by Xilinx and must be used           --
--     solely for design, simulation, implementation and creation of          --
--     design files limited to Xilinx devices or technologies. Use            --
--     with non-Xilinx devices or technologies is expressly prohibited        --
--     and immediately terminates your license.                               --
--                                                                            --
--     XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS"          --
--     SOLELY FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR                --
--     XILINX DEVICES.  BY PROVIDING THIS DESIGN, CODE, OR INFORMATION        --
--     AS ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE, APPLICATION            --
--     OR STANDARD, XILINX IS MAKING NO REPRESENTATION THAT THIS              --
--     IMPLEMENTATION IS FREE FROM ANY CLAIMS OF INFRINGEMENT,                --
--     AND YOU ARE RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY REQUIRE       --
--     FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY DISCLAIMS ANY               --
--     WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE                --
--     IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR         --
--     REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF        --
--     INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS        --
--     FOR A PARTICULAR PURPOSE.                                              --
--                                                                            --
--     Xilinx products are not intended for use in life support               --
--     appliances, devices, or systems. Use in such applications are          --
--     expressly prohibited.                                                  --
--                                                                            --
--     (c) Copyright 1995-2006 Xilinx, Inc.                                   --
--     All rights reserved.                                                   --
--------------------------------------------------------------------------------

-- synthesis translate_off
LIBRARY std, ieee;
USE std.standard.ALL;
USE ieee.std_logic_1164.ALL;

LIBRARY unisim;
USE unisim.vcomponents.ALL;


LIBRARY XilinxCoreLib;
USE XilinxCoreLib.c_addsub_v5_0_comp.ALL;
USE XilinxCoreLib.c_da_fir_v7_0_comp.ALL;
USE XilinxCoreLib.c_mux_bus_v5_0_comp.ALL;
USE XilinxCoreLib.c_counter_binary_v5_0_comp.ALL;
USE XilinxCoreLib.c_cic_v3_0_comp.ALL;
USE XilinxCoreLib.c_reg_fd_v5_0_comp.ALL;
USE XilinxCoreLib.c_dds_v4_1_comp.ALL;
USE XilinxCoreLib.c_shift_ram_v5_0_comp.ALL;
USE XilinxCoreLib.mult_gen_v5_0_comp.ALL;
USE XilinxCoreLib.c_gate_bit_v5_0_comp.ALL;

ENTITY myddc IS
   PORT (
      DIN : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
      ND : IN STD_LOGIC;
      CLK : IN STD_LOGIC;
      ADDR : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      LD_DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      WE : IN STD_LOGIC;
      SEL : IN STD_LOGIC;
      RDY : OUT STD_LOGIC;
      RFD : OUT STD_LOGIC;
      DOUT_I : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
      DOUT_Q : OUT STD_LOGIC_VECTOR(29 DOWNTO 0)   
);
END myddc;

ARCHITECTURE xilinx OF myddc IS 

-- Signals for connecting to instantiations
   SIGNAL BU4_I0 : STD_LOGIC;
   SIGNAL BU4_I1 : STD_LOGIC;
   SIGNAL BU4_I2 : STD_LOGIC;
   SIGNAL BU4_I3 : STD_LOGIC;
   SIGNAL BU4_O : STD_LOGIC;
   SIGNAL BU8_I0 : STD_LOGIC;
   SIGNAL BU8_I1 : STD_LOGIC;
   SIGNAL BU8_I2 : STD_LOGIC;
   SIGNAL BU8_I3 : STD_LOGIC;
   SIGNAL BU8_O : STD_LOGIC;
   SIGNAL BU10_I0 : STD_LOGIC;
   SIGNAL BU10_I1 : STD_LOGIC;
   SIGNAL BU10_I2 : STD_LOGIC;
   SIGNAL BU10_I3 : STD_LOGIC;
   SIGNAL BU10_O : STD_LOGIC;
   SIGNAL BU1292_D : STD_LOGIC;
   SIGNAL BU1292_C : STD_LOGIC;
   SIGNAL BU1292_CE : STD_LOGIC;
   SIGNAL BU1292_Q : STD_LOGIC;
   SIGNAL BU14_D : STD_LOGIC;
   SIGNAL BU14_CE : STD_LOGIC;
   SIGNAL BU14_CLK : STD_LOGIC;
   SIGNAL BU14_A0 : STD_LOGIC;
   SIGNAL BU14_A1 : STD_LOGIC;
   SIGNAL BU14_A2 : STD_LOGIC;
   SIGNAL BU14_A3 : STD_LOGIC;
   SIGNAL BU14_Q : STD_LOGIC;
   SIGNAL BU16_D : STD_LOGIC;
   SIGNAL BU16_C : STD_LOGIC;
   SIGNAL BU16_CE : STD_LOGIC;
   SIGNAL BU16_Q : STD_LOGIC;
   SIGNAL BU17_D : STD_LOGIC;
   SIGNAL BU17_CE : STD_LOGIC;
   SIGNAL BU17_CLK : STD_LOGIC;
   SIGNAL BU17_A0 : STD_LOGIC;
   SIGNAL BU17_A1 : STD_LOGIC;
   SIGNAL BU17_A2 : STD_LOGIC;
   SIGNAL BU17_A3 : STD_LOGIC;
   SIGNAL BU17_Q : STD_LOGIC;
   SIGNAL BU19_D : STD_LOGIC;
   SIGNAL BU19_C : STD_LOGIC;
   SIGNAL BU19_CE : STD_LOGIC;
   SIGNAL BU19_Q : STD_LOGIC;
   SIGNAL BU20_D : STD_LOGIC;
   SIGNAL BU20_CE : STD_LOGIC;
   SIGNAL BU20_CLK : STD_LOGIC;
   SIGNAL BU20_A0 : STD_LOGIC;
   SIGNAL BU20_A1 : STD_LOGIC;
   SIGNAL BU20_A2 : STD_LOGIC;
   SIGNAL BU20_A3 : STD_LOGIC;
   SIGNAL BU20_Q : STD_LOGIC;
   SIGNAL BU22_D : STD_LOGIC;
   SIGNAL BU22_C : STD_LOGIC;
   SIGNAL BU22_CE : STD_LOGIC;
   SIGNAL BU22_Q : STD_LOGIC;
   SIGNAL BU23_D : STD_LOGIC;
   SIGNAL BU23_CE : STD_LOGIC;
   SIGNAL BU23_CLK : STD_LOGIC;
   SIGNAL BU23_A0 : STD_LOGIC;
   SIGNAL BU23_A1 : STD_LOGIC;
   SIGNAL BU23_A2 : STD_LOGIC;
   SIGNAL BU23_A3 : STD_LOGIC;
   SIGNAL BU23_Q : STD_LOGIC;
   SIGNAL BU25_D : STD_LOGIC;
   SIGNAL BU25_C : STD_LOGIC;
   SIGNAL BU25_CE : STD_LOGIC;
   SIGNAL BU25_Q : STD_LOGIC;
   SIGNAL BU26_D : STD_LOGIC;
   SIGNAL BU26_CE : STD_LOGIC;
   SIGNAL BU26_CLK : STD_LOGIC;
   SIGNAL BU26_A0 : STD_LOGIC;
   SIGNAL BU26_A1 : STD_LOGIC;
   SIGNAL BU26_A2 : STD_LOGIC;
   SIGNAL BU26_A3 : STD_LOGIC;
   SIGNAL BU26_Q : STD_LOGIC;
   SIGNAL BU28_D : STD_LOGIC;
   SIGNAL BU28_C : STD_LOGIC;
   SIGNAL BU28_CE : STD_LOGIC;
   SIGNAL BU28_Q : STD_LOGIC;
   SIGNAL BU29_D : STD_LOGIC;
   SIGNAL BU29_CE : STD_LOGIC;
   SIGNAL BU29_CLK : STD_LOGIC;
   SIGNAL BU29_A0 : STD_LOGIC;
   SIGNAL BU29_A1 : STD_LOGIC;
   SIGNAL BU29_A2 : STD_LOGIC;
   SIGNAL BU29_A3 : STD_LOGIC;
   SIGNAL BU29_Q : STD_LOGIC;
   SIGNAL BU31_D : STD_LOGIC;
   SIGNAL BU31_C : STD_LOGIC;
   SIGNAL BU31_CE : STD_LOGIC;
   SIGNAL BU31_Q : STD_LOGIC;
   SIGNAL BU32_D : STD_LOGIC;
   SIGNAL BU32_CE : STD_LOGIC;
   SIGNAL BU32_CLK : STD_LOGIC;
   SIGNAL BU32_A0 : STD_LOGIC;
   SIGNAL BU32_A1 : STD_LOGIC;
   SIGNAL BU32_A2 : STD_LOGIC;
   SIGNAL BU32_A3 : STD_LOGIC;
   SIGNAL BU32_Q : STD_LOGIC;
   SIGNAL BU34_D : STD_LOGIC;
   SIGNAL BU34_C : STD_LOGIC;
   SIGNAL BU34_CE : STD_LOGIC;
   SIGNAL BU34_Q : STD_LOGIC;
   SIGNAL BU35_D : STD_LOGIC;
   SIGNAL BU35_CE : STD_LOGIC;
   SIGNAL BU35_CLK : STD_LOGIC;
   SIGNAL BU35_A0 : STD_LOGIC;
   SIGNAL BU35_A1 : STD_LOGIC;
   SIGNAL BU35_A2 : STD_LOGIC;
   SIGNAL BU35_A3 : STD_LOGIC;
   SIGNAL BU35_Q : STD_LOGIC;
   SIGNAL BU37_D : STD_LOGIC;
   SIGNAL BU37_C : STD_LOGIC;
   SIGNAL BU37_CE : STD_LOGIC;
   SIGNAL BU37_Q : STD_LOGIC;
   SIGNAL BU38_D : STD_LOGIC;
   SIGNAL BU38_CE : STD_LOGIC;
   SIGNAL BU38_CLK : STD_LOGIC;
   SIGNAL BU38_A0 : STD_LOGIC;
   SIGNAL BU38_A1 : STD_LOGIC;
   SIGNAL BU38_A2 : STD_LOGIC;
   SIGNAL BU38_A3 : STD_LOGIC;
   SIGNAL BU38_Q : STD_LOGIC;
   SIGNAL BU40_D : STD_LOGIC;
   SIGNAL BU40_C : STD_LOGIC;
   SIGNAL BU40_CE : STD_LOGIC;
   SIGNAL BU40_Q : STD_LOGIC;
   SIGNAL BU41_D : STD_LOGIC;
   SIGNAL BU41_CE : STD_LOGIC;
   SIGNAL BU41_CLK : STD_LOGIC;
   SIGNAL BU41_A0 : STD_LOGIC;
   SIGNAL BU41_A1 : STD_LOGIC;
   SIGNAL BU41_A2 : STD_LOGIC;
   SIGNAL BU41_A3 : STD_LOGIC;
   SIGNAL BU41_Q : STD_LOGIC;
   SIGNAL BU43_D : STD_LOGIC;
   SIGNAL BU43_C : STD_LOGIC;
   SIGNAL BU43_CE : STD_LOGIC;
   SIGNAL BU43_Q : STD_LOGIC;
   SIGNAL BU44_D : STD_LOGIC;
   SIGNAL BU44_CE : STD_LOGIC;
   SIGNAL BU44_CLK : STD_LOGIC;
   SIGNAL BU44_A0 : STD_LOGIC;
   SIGNAL BU44_A1 : STD_LOGIC;
   SIGNAL BU44_A2 : STD_LOGIC;
   SIGNAL BU44_A3 : STD_LOGIC;
   SIGNAL BU44_Q : STD_LOGIC;
   SIGNAL BU46_D : STD_LOGIC;
   SIGNAL BU46_C : STD_LOGIC;
   SIGNAL BU46_CE : STD_LOGIC;
   SIGNAL BU46_Q : STD_LOGIC;
   SIGNAL BU47_D : STD_LOGIC;
   SIGNAL BU47_CE : STD_LOGIC;
   SIGNAL BU47_CLK : STD_LOGIC;
   SIGNAL BU47_A0 : STD_LOGIC;
   SIGNAL BU47_A1 : STD_LOGIC;
   SIGNAL BU47_A2 : STD_LOGIC;
   SIGNAL BU47_A3 : STD_LOGIC;
   SIGNAL BU47_Q : STD_LOGIC;
   SIGNAL BU49_D : STD_LOGIC;
   SIGNAL BU49_C : STD_LOGIC;
   SIGNAL BU49_CE : STD_LOGIC;
   SIGNAL BU49_Q : STD_LOGIC;
   SIGNAL BU50_D : STD_LOGIC;
   SIGNAL BU50_CE : STD_LOGIC;
   SIGNAL BU50_CLK : STD_LOGIC;
   SIGNAL BU50_A0 : STD_LOGIC;
   SIGNAL BU50_A1 : STD_LOGIC;
   SIGNAL BU50_A2 : STD_LOGIC;
   SIGNAL BU50_A3 : STD_LOGIC;
   SIGNAL BU50_Q : STD_LOGIC;
   SIGNAL BU52_D : STD_LOGIC;
   SIGNAL BU52_C : STD_LOGIC;
   SIGNAL BU52_CE : STD_LOGIC;
   SIGNAL BU52_Q : STD_LOGIC;
   SIGNAL BU53_D : STD_LOGIC;
   SIGNAL BU53_CE : STD_LOGIC;
   SIGNAL BU53_CLK : STD_LOGIC;
   SIGNAL BU53_A0 : STD_LOGIC;
   SIGNAL BU53_A1 : STD_LOGIC;
   SIGNAL BU53_A2 : STD_LOGIC;
   SIGNAL BU53_A3 : STD_LOGIC;
   SIGNAL BU53_Q : STD_LOGIC;
   SIGNAL BU55_D : STD_LOGIC;
   SIGNAL BU55_C : STD_LOGIC;
   SIGNAL BU55_CE : STD_LOGIC;
   SIGNAL BU55_Q : STD_LOGIC;
   SIGNAL BU57_DATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
   SIGNAL BU57_WE : STD_LOGIC;
   SIGNAL BU57_CLK : STD_LOGIC;
   SIGNAL BU57_CE : STD_LOGIC;
   SIGNAL BU57_RDY : STD_LOGIC;
   SIGNAL BU57_SINE : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU57_COSINE : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1294_I0 : STD_LOGIC;
   SIGNAL BU1294_I1 : STD_LOGIC;
   SIGNAL BU1294_I2 : STD_LOGIC;
   SIGNAL BU1294_I3 : STD_LOGIC;
   SIGNAL BU1294_O : STD_LOGIC;
   SIGNAL BU1296_clk : STD_LOGIC;
   SIGNAL BU1296_a : STD_LOGIC_VECTOR(13 DOWNTO 0);
   SIGNAL BU1296_b : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1296_o : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1296_q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1296_a_signed : STD_LOGIC;
   SIGNAL BU1296_loadb : STD_LOGIC;
   SIGNAL BU1296_load_done : STD_LOGIC;
   SIGNAL BU1296_swapb : STD_LOGIC;
   SIGNAL BU1296_ce : STD_LOGIC;
   SIGNAL BU1296_aclr : STD_LOGIC;
   SIGNAL BU1296_sclr : STD_LOGIC;
   SIGNAL BU1296_rfd : STD_LOGIC;
   SIGNAL BU1296_nd : STD_LOGIC;
   SIGNAL BU1296_rdy : STD_LOGIC;
   SIGNAL BU1517_I : STD_LOGIC_VECTOR(4 DOWNTO 0);
   SIGNAL BU1517_O : STD_LOGIC;
   SIGNAL BU1526_I0 : STD_LOGIC;
   SIGNAL BU1526_I1 : STD_LOGIC;
   SIGNAL BU1526_I2 : STD_LOGIC;
   SIGNAL BU1526_I3 : STD_LOGIC;
   SIGNAL BU1526_O : STD_LOGIC;
   SIGNAL BU1527_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU1527_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1527_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU1628_I0 : STD_LOGIC;
   SIGNAL BU1628_I1 : STD_LOGIC;
   SIGNAL BU1628_I2 : STD_LOGIC;
   SIGNAL BU1628_I3 : STD_LOGIC;
   SIGNAL BU1628_O : STD_LOGIC;
   SIGNAL BU1630_I0 : STD_LOGIC;
   SIGNAL BU1630_I1 : STD_LOGIC;
   SIGNAL BU1630_I2 : STD_LOGIC;
   SIGNAL BU1630_I3 : STD_LOGIC;
   SIGNAL BU1630_O : STD_LOGIC;
   SIGNAL BU1631_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU1631_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU1631_CLK : STD_LOGIC;
   SIGNAL BU1631_SCLR : STD_LOGIC;
   SIGNAL BU1631_SSET : STD_LOGIC;
   SIGNAL BU1724_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1724_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1724_CLK : STD_LOGIC;
   SIGNAL BU1724_SCLR : STD_LOGIC;
   SIGNAL BU1724_SSET : STD_LOGIC;
   SIGNAL BU1729_CLK : STD_LOGIC;
   SIGNAL BU1729_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1729_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1734_clk : STD_LOGIC;
   SIGNAL BU1734_a : STD_LOGIC_VECTOR(13 DOWNTO 0);
   SIGNAL BU1734_b : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1734_o : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1734_q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1734_a_signed : STD_LOGIC;
   SIGNAL BU1734_loadb : STD_LOGIC;
   SIGNAL BU1734_load_done : STD_LOGIC;
   SIGNAL BU1734_swapb : STD_LOGIC;
   SIGNAL BU1734_ce : STD_LOGIC;
   SIGNAL BU1734_aclr : STD_LOGIC;
   SIGNAL BU1734_sclr : STD_LOGIC;
   SIGNAL BU1734_rfd : STD_LOGIC;
   SIGNAL BU1734_nd : STD_LOGIC;
   SIGNAL BU1734_rdy : STD_LOGIC;
   SIGNAL BU1955_I : STD_LOGIC_VECTOR(4 DOWNTO 0);
   SIGNAL BU1955_O : STD_LOGIC;
   SIGNAL BU1964_I0 : STD_LOGIC;
   SIGNAL BU1964_I1 : STD_LOGIC;
   SIGNAL BU1964_I2 : STD_LOGIC;
   SIGNAL BU1964_I3 : STD_LOGIC;
   SIGNAL BU1964_O : STD_LOGIC;
   SIGNAL BU1965_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU1965_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1965_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU2066_I0 : STD_LOGIC;
   SIGNAL BU2066_I1 : STD_LOGIC;
   SIGNAL BU2066_I2 : STD_LOGIC;
   SIGNAL BU2066_I3 : STD_LOGIC;
   SIGNAL BU2066_O : STD_LOGIC;
   SIGNAL BU2068_I0 : STD_LOGIC;
   SIGNAL BU2068_I1 : STD_LOGIC;
   SIGNAL BU2068_I2 : STD_LOGIC;
   SIGNAL BU2068_I3 : STD_LOGIC;
   SIGNAL BU2068_O : STD_LOGIC;
   SIGNAL BU2069_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2069_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2069_CLK : STD_LOGIC;
   SIGNAL BU2069_SCLR : STD_LOGIC;
   SIGNAL BU2069_SSET : STD_LOGIC;
   SIGNAL BU2162_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2162_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2162_CLK : STD_LOGIC;
   SIGNAL BU2162_SCLR : STD_LOGIC;
   SIGNAL BU2162_SSET : STD_LOGIC;
   SIGNAL BU2457_D : STD_LOGIC;
   SIGNAL BU2457_C : STD_LOGIC;
   SIGNAL BU2457_CE : STD_LOGIC;
   SIGNAL BU2457_Q : STD_LOGIC;
   SIGNAL BU2461_I : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2461_O : STD_LOGIC;
   SIGNAL BU2489_I0 : STD_LOGIC;
   SIGNAL BU2489_I1 : STD_LOGIC;
   SIGNAL BU2489_I2 : STD_LOGIC;
   SIGNAL BU2489_I3 : STD_LOGIC;
   SIGNAL BU2489_O : STD_LOGIC;
   SIGNAL BU2490_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2490_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2490_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU2591_I0 : STD_LOGIC;
   SIGNAL BU2591_I1 : STD_LOGIC;
   SIGNAL BU2591_I2 : STD_LOGIC;
   SIGNAL BU2591_I3 : STD_LOGIC;
   SIGNAL BU2591_O : STD_LOGIC;
   SIGNAL BU2593_I0 : STD_LOGIC;
   SIGNAL BU2593_I1 : STD_LOGIC;
   SIGNAL BU2593_I2 : STD_LOGIC;
   SIGNAL BU2593_I3 : STD_LOGIC;
   SIGNAL BU2593_O : STD_LOGIC;
   SIGNAL BU2594_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2594_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2594_CLK : STD_LOGIC;
   SIGNAL BU2594_SCLR : STD_LOGIC;
   SIGNAL BU2594_SSET : STD_LOGIC;
   SIGNAL BU2687_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2687_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2687_CLK : STD_LOGIC;
   SIGNAL BU2687_SCLR : STD_LOGIC;
   SIGNAL BU2687_SSET : STD_LOGIC;
   SIGNAL BU7487_I : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU7487_O : STD_LOGIC;
   SIGNAL BU7515_I0 : STD_LOGIC;
   SIGNAL BU7515_I1 : STD_LOGIC;
   SIGNAL BU7515_I2 : STD_LOGIC;
   SIGNAL BU7515_I3 : STD_LOGIC;
   SIGNAL BU7515_O : STD_LOGIC;
   SIGNAL BU7516_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU7516_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU7516_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU7617_I0 : STD_LOGIC;
   SIGNAL BU7617_I1 : STD_LOGIC;
   SIGNAL BU7617_I2 : STD_LOGIC;
   SIGNAL BU7617_I3 : STD_LOGIC;
   SIGNAL BU7617_O : STD_LOGIC;
   SIGNAL BU7619_I0 : STD_LOGIC;
   SIGNAL BU7619_I1 : STD_LOGIC;
   SIGNAL BU7619_I2 : STD_LOGIC;
   SIGNAL BU7619_I3 : STD_LOGIC;
   SIGNAL BU7619_O : STD_LOGIC;
   SIGNAL BU7620_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU7620_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU7620_CLK : STD_LOGIC;
   SIGNAL BU7620_SCLR : STD_LOGIC;
   SIGNAL BU7620_SSET : STD_LOGIC;
   SIGNAL BU7713_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU7713_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU7713_CLK : STD_LOGIC;
   SIGNAL BU7713_SCLR : STD_LOGIC;
   SIGNAL BU7713_SSET : STD_LOGIC;
   SIGNAL BU2173_D : STD_LOGIC;
   SIGNAL BU2173_C : STD_LOGIC;
   SIGNAL BU2173_CE : STD_LOGIC;
   SIGNAL BU2173_Q : STD_LOGIC;
   SIGNAL BU2175_D : STD_LOGIC;
   SIGNAL BU2175_C : STD_LOGIC;
   SIGNAL BU2175_CE : STD_LOGIC;
   SIGNAL BU2175_Q : STD_LOGIC;
   SIGNAL BU2177_D : STD_LOGIC;
   SIGNAL BU2177_C : STD_LOGIC;
   SIGNAL BU2177_CE : STD_LOGIC;
   SIGNAL BU2177_Q : STD_LOGIC;
   SIGNAL BU2179_D : STD_LOGIC;
   SIGNAL BU2179_C : STD_LOGIC;
   SIGNAL BU2179_CE : STD_LOGIC;
   SIGNAL BU2179_Q : STD_LOGIC;
   SIGNAL BU2181_D : STD_LOGIC;
   SIGNAL BU2181_C : STD_LOGIC;
   SIGNAL BU2181_CE : STD_LOGIC;
   SIGNAL BU2181_Q : STD_LOGIC;
   SIGNAL BU2183_D : STD_LOGIC;
   SIGNAL BU2183_C : STD_LOGIC;
   SIGNAL BU2183_CE : STD_LOGIC;
   SIGNAL BU2183_Q : STD_LOGIC;
   SIGNAL BU2185_D : STD_LOGIC;
   SIGNAL BU2185_C : STD_LOGIC;
   SIGNAL BU2185_CE : STD_LOGIC;
   SIGNAL BU2185_Q : STD_LOGIC;
   SIGNAL BU2187_D : STD_LOGIC;
   SIGNAL BU2187_C : STD_LOGIC;
   SIGNAL BU2187_CE : STD_LOGIC;
   SIGNAL BU2187_Q : STD_LOGIC;
   SIGNAL BU2189_D : STD_LOGIC;
   SIGNAL BU2189_C : STD_LOGIC;
   SIGNAL BU2189_CE : STD_LOGIC;
   SIGNAL BU2189_Q : STD_LOGIC;
   SIGNAL BU2191_D : STD_LOGIC;
   SIGNAL BU2191_C : STD_LOGIC;
   SIGNAL BU2191_CE : STD_LOGIC;
   SIGNAL BU2191_Q : STD_LOGIC;
   SIGNAL BU2193_D : STD_LOGIC;
   SIGNAL BU2193_C : STD_LOGIC;
   SIGNAL BU2193_CE : STD_LOGIC;
   SIGNAL BU2193_Q : STD_LOGIC;
   SIGNAL BU2195_D : STD_LOGIC;
   SIGNAL BU2195_C : STD_LOGIC;
   SIGNAL BU2195_CE : STD_LOGIC;
   SIGNAL BU2195_Q : STD_LOGIC;
   SIGNAL BU2197_D : STD_LOGIC;
   SIGNAL BU2197_C : STD_LOGIC;
   SIGNAL BU2197_CE : STD_LOGIC;
   SIGNAL BU2197_Q : STD_LOGIC;
   SIGNAL BU2199_D : STD_LOGIC;
   SIGNAL BU2199_C : STD_LOGIC;
   SIGNAL BU2199_CE : STD_LOGIC;
   SIGNAL BU2199_Q : STD_LOGIC;
   SIGNAL BU2201_D : STD_LOGIC;
   SIGNAL BU2201_C : STD_LOGIC;
   SIGNAL BU2201_CE : STD_LOGIC;
   SIGNAL BU2201_Q : STD_LOGIC;
   SIGNAL BU2203_D : STD_LOGIC;
   SIGNAL BU2203_C : STD_LOGIC;
   SIGNAL BU2203_CE : STD_LOGIC;
   SIGNAL BU2203_Q : STD_LOGIC;
   SIGNAL BU2205_D : STD_LOGIC;
   SIGNAL BU2205_C : STD_LOGIC;
   SIGNAL BU2205_CE : STD_LOGIC;
   SIGNAL BU2205_Q : STD_LOGIC;
   SIGNAL BU2207_D : STD_LOGIC;
   SIGNAL BU2207_C : STD_LOGIC;
   SIGNAL BU2207_CE : STD_LOGIC;
   SIGNAL BU2207_Q : STD_LOGIC;
   SIGNAL BU2209_D : STD_LOGIC;
   SIGNAL BU2209_C : STD_LOGIC;
   SIGNAL BU2209_CE : STD_LOGIC;
   SIGNAL BU2209_Q : STD_LOGIC;
   SIGNAL BU2211_D : STD_LOGIC;
   SIGNAL BU2211_C : STD_LOGIC;
   SIGNAL BU2211_CE : STD_LOGIC;
   SIGNAL BU2211_Q : STD_LOGIC;
   SIGNAL BU2213_D : STD_LOGIC;
   SIGNAL BU2213_C : STD_LOGIC;
   SIGNAL BU2213_CE : STD_LOGIC;
   SIGNAL BU2213_Q : STD_LOGIC;
   SIGNAL BU2215_D : STD_LOGIC;
   SIGNAL BU2215_C : STD_LOGIC;
   SIGNAL BU2215_CE : STD_LOGIC;
   SIGNAL BU2215_Q : STD_LOGIC;
   SIGNAL BU2217_D : STD_LOGIC;
   SIGNAL BU2217_C : STD_LOGIC;
   SIGNAL BU2217_CE : STD_LOGIC;
   SIGNAL BU2217_Q : STD_LOGIC;
   SIGNAL BU2219_D : STD_LOGIC;
   SIGNAL BU2219_C : STD_LOGIC;
   SIGNAL BU2219_CE : STD_LOGIC;
   SIGNAL BU2219_Q : STD_LOGIC;
   SIGNAL BU2220_MA : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_MB : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_S : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2220_Q : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_CLK : STD_LOGIC;
   SIGNAL BU2448_D : STD_LOGIC;
   SIGNAL BU2448_C : STD_LOGIC;
   SIGNAL BU2448_CE : STD_LOGIC;
   SIGNAL BU2448_Q : STD_LOGIC;
   SIGNAL BU2452_I0 : STD_LOGIC;
   SIGNAL BU2452_I1 : STD_LOGIC;
   SIGNAL BU2452_I2 : STD_LOGIC;
   SIGNAL BU2452_I3 : STD_LOGIC;
   SIGNAL BU2452_O : STD_LOGIC;
   SIGNAL BU2453_D : STD_LOGIC;
   SIGNAL BU2453_C : STD_LOGIC;
   SIGNAL BU2453_CE : STD_LOGIC;
   SIGNAL BU2453_Q : STD_LOGIC;
   SIGNAL BU2692_DIN : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2692_ND : STD_LOGIC;
   SIGNAL BU2692_RFD : STD_LOGIC;
   SIGNAL BU2692_CLK : STD_LOGIC;
   SIGNAL BU2692_DOUT : STD_LOGIC_VECTOR(46 DOWNTO 0);
   SIGNAL BU2692_RDY : STD_LOGIC;
   SIGNAL BU7718_DIN : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU7718_ND : STD_LOGIC;
   SIGNAL BU7718_RFD : STD_LOGIC;
   SIGNAL BU7718_CLK : STD_LOGIC;
   SIGNAL BU7718_DOUT : STD_LOGIC_VECTOR(46 DOWNTO 0);
   SIGNAL BU7718_RDY : STD_LOGIC;
   SIGNAL BU12513_I0 : STD_LOGIC;
   SIGNAL BU12513_I1 : STD_LOGIC;
   SIGNAL BU12513_I2 : STD_LOGIC;
   SIGNAL BU12513_I3 : STD_LOGIC;
   SIGNAL BU12513_O : STD_LOGIC;
   SIGNAL BU12518_I0 : STD_LOGIC;
   SIGNAL BU12518_I1 : STD_LOGIC;
   SIGNAL BU12518_I2 : STD_LOGIC;
   SIGNAL BU12518_I3 : STD_LOGIC;
   SIGNAL BU12518_O : STD_LOGIC;
   SIGNAL BU12524_D : STD_LOGIC;
   SIGNAL BU12524_CE : STD_LOGIC;
   SIGNAL BU12524_CLK : STD_LOGIC;
   SIGNAL BU12524_A0 : STD_LOGIC;
   SIGNAL BU12524_A1 : STD_LOGIC;
   SIGNAL BU12524_A2 : STD_LOGIC;
   SIGNAL BU12524_A3 : STD_LOGIC;
   SIGNAL BU12524_Q : STD_LOGIC;
   SIGNAL BU12525_D : STD_LOGIC;
   SIGNAL BU12525_CE : STD_LOGIC;
   SIGNAL BU12525_CLK : STD_LOGIC;
   SIGNAL BU12525_A0 : STD_LOGIC;
   SIGNAL BU12525_A1 : STD_LOGIC;
   SIGNAL BU12525_A2 : STD_LOGIC;
   SIGNAL BU12525_A3 : STD_LOGIC;
   SIGNAL BU12525_Q : STD_LOGIC;
   SIGNAL BU12526_D : STD_LOGIC;
   SIGNAL BU12526_CE : STD_LOGIC;
   SIGNAL BU12526_CLK : STD_LOGIC;
   SIGNAL BU12526_A0 : STD_LOGIC;
   SIGNAL BU12526_A1 : STD_LOGIC;
   SIGNAL BU12526_A2 : STD_LOGIC;
   SIGNAL BU12526_A3 : STD_LOGIC;
   SIGNAL BU12526_Q : STD_LOGIC;
   SIGNAL BU12527_D : STD_LOGIC;
   SIGNAL BU12527_CE : STD_LOGIC;
   SIGNAL BU12527_CLK : STD_LOGIC;
   SIGNAL BU12527_A0 : STD_LOGIC;
   SIGNAL BU12527_A1 : STD_LOGIC;
   SIGNAL BU12527_A2 : STD_LOGIC;
   SIGNAL BU12527_A3 : STD_LOGIC;
   SIGNAL BU12527_Q : STD_LOGIC;
   SIGNAL BU12528_D : STD_LOGIC;
   SIGNAL BU12528_CE : STD_LOGIC;
   SIGNAL BU12528_CLK : STD_LOGIC;
   SIGNAL BU12528_A0 : STD_LOGIC;
   SIGNAL BU12528_A1 : STD_LOGIC;
   SIGNAL BU12528_A2 : STD_LOGIC;
   SIGNAL BU12528_A3 : STD_LOGIC;
   SIGNAL BU12528_Q : STD_LOGIC;
   SIGNAL BU12529_D : STD_LOGIC;
   SIGNAL BU12529_CE : STD_LOGIC;
   SIGNAL BU12529_CLK : STD_LOGIC;
   SIGNAL BU12529_A0 : STD_LOGIC;
   SIGNAL BU12529_A1 : STD_LOGIC;
   SIGNAL BU12529_A2 : STD_LOGIC;
   SIGNAL BU12529_A3 : STD_LOGIC;
   SIGNAL BU12529_Q : STD_LOGIC;
   SIGNAL BU12530_D : STD_LOGIC;
   SIGNAL BU12530_CE : STD_LOGIC;
   SIGNAL BU12530_CLK : STD_LOGIC;
   SIGNAL BU12530_A0 : STD_LOGIC;
   SIGNAL BU12530_A1 : STD_LOGIC;
   SIGNAL BU12530_A2 : STD_LOGIC;
   SIGNAL BU12530_A3 : STD_LOGIC;
   SIGNAL BU12530_Q : STD_LOGIC;
   SIGNAL BU12531_D : STD_LOGIC;
   SIGNAL BU12531_CE : STD_LOGIC;
   SIGNAL BU12531_CLK : STD_LOGIC;
   SIGNAL BU12531_A0 : STD_LOGIC;
   SIGNAL BU12531_A1 : STD_LOGIC;
   SIGNAL BU12531_A2 : STD_LOGIC;
   SIGNAL BU12531_A3 : STD_LOGIC;
   SIGNAL BU12531_Q : STD_LOGIC;
   SIGNAL BU12532_D : STD_LOGIC;
   SIGNAL BU12532_CE : STD_LOGIC;
   SIGNAL BU12532_CLK : STD_LOGIC;
   SIGNAL BU12532_A0 : STD_LOGIC;
   SIGNAL BU12532_A1 : STD_LOGIC;
   SIGNAL BU12532_A2 : STD_LOGIC;
   SIGNAL BU12532_A3 : STD_LOGIC;
   SIGNAL BU12532_Q : STD_LOGIC;
   SIGNAL BU12533_D : STD_LOGIC;
   SIGNAL BU12533_CE : STD_LOGIC;
   SIGNAL BU12533_CLK : STD_LOGIC;
   SIGNAL BU12533_A0 : STD_LOGIC;
   SIGNAL BU12533_A1 : STD_LOGIC;
   SIGNAL BU12533_A2 : STD_LOGIC;
   SIGNAL BU12533_A3 : STD_LOGIC;
   SIGNAL BU12533_Q : STD_LOGIC;
   SIGNAL BU12534_D : STD_LOGIC;
   SIGNAL BU12534_CE : STD_LOGIC;
   SIGNAL BU12534_CLK : STD_LOGIC;
   SIGNAL BU12534_A0 : STD_LOGIC;
   SIGNAL BU12534_A1 : STD_LOGIC;
   SIGNAL BU12534_A2 : STD_LOGIC;
   SIGNAL BU12534_A3 : STD_LOGIC;
   SIGNAL BU12534_Q : STD_LOGIC;
   SIGNAL BU12535_D : STD_LOGIC;
   SIGNAL BU12535_CE : STD_LOGIC;
   SIGNAL BU12535_CLK : STD_LOGIC;
   SIGNAL BU12535_A0 : STD_LOGIC;
   SIGNAL BU12535_A1 : STD_LOGIC;
   SIGNAL BU12535_A2 : STD_LOGIC;
   SIGNAL BU12535_A3 : STD_LOGIC;
   SIGNAL BU12535_Q : STD_LOGIC;
   SIGNAL BU12536_D : STD_LOGIC;
   SIGNAL BU12536_CE : STD_LOGIC;
   SIGNAL BU12536_CLK : STD_LOGIC;
   SIGNAL BU12536_A0 : STD_LOGIC;
   SIGNAL BU12536_A1 : STD_LOGIC;
   SIGNAL BU12536_A2 : STD_LOGIC;
   SIGNAL BU12536_A3 : STD_LOGIC;
   SIGNAL BU12536_Q : STD_LOGIC;
   SIGNAL BU12537_D : STD_LOGIC;
   SIGNAL BU12537_CE : STD_LOGIC;
   SIGNAL BU12537_CLK : STD_LOGIC;
   SIGNAL BU12537_A0 : STD_LOGIC;
   SIGNAL BU12537_A1 : STD_LOGIC;
   SIGNAL BU12537_A2 : STD_LOGIC;
   SIGNAL BU12537_A3 : STD_LOGIC;
   SIGNAL BU12537_Q : STD_LOGIC;
   SIGNAL BU12538_D : STD_LOGIC;
   SIGNAL BU12538_CE : STD_LOGIC;
   SIGNAL BU12538_CLK : STD_LOGIC;
   SIGNAL BU12538_A0 : STD_LOGIC;
   SIGNAL BU12538_A1 : STD_LOGIC;
   SIGNAL BU12538_A2 : STD_LOGIC;
   SIGNAL BU12538_A3 : STD_LOGIC;
   SIGNAL BU12538_Q : STD_LOGIC;
   SIGNAL BU12539_D : STD_LOGIC;
   SIGNAL BU12539_CE : STD_LOGIC;
   SIGNAL BU12539_CLK : STD_LOGIC;
   SIGNAL BU12539_A0 : STD_LOGIC;
   SIGNAL BU12539_A1 : STD_LOGIC;
   SIGNAL BU12539_A2 : STD_LOGIC;
   SIGNAL BU12539_A3 : STD_LOGIC;
   SIGNAL BU12539_Q : STD_LOGIC;
   SIGNAL BU12540_D : STD_LOGIC;
   SIGNAL BU12540_CE : STD_LOGIC;
   SIGNAL BU12540_CLK : STD_LOGIC;
   SIGNAL BU12540_A0 : STD_LOGIC;
   SIGNAL BU12540_A1 : STD_LOGIC;
   SIGNAL BU12540_A2 : STD_LOGIC;
   SIGNAL BU12540_A3 : STD_LOGIC;
   SIGNAL BU12540_Q : STD_LOGIC;
   SIGNAL BU12541_D : STD_LOGIC;
   SIGNAL BU12541_CE : STD_LOGIC;
   SIGNAL BU12541_CLK : STD_LOGIC;
   SIGNAL BU12541_A0 : STD_LOGIC;
   SIGNAL BU12541_A1 : STD_LOGIC;
   SIGNAL BU12541_A2 : STD_LOGIC;
   SIGNAL BU12541_A3 : STD_LOGIC;
   SIGNAL BU12541_Q : STD_LOGIC;
   SIGNAL BU12542_D : STD_LOGIC;
   SIGNAL BU12542_CE : STD_LOGIC;
   SIGNAL BU12542_CLK : STD_LOGIC;
   SIGNAL BU12542_A0 : STD_LOGIC;
   SIGNAL BU12542_A1 : STD_LOGIC;
   SIGNAL BU12542_A2 : STD_LOGIC;
   SIGNAL BU12542_A3 : STD_LOGIC;
   SIGNAL BU12542_Q : STD_LOGIC;
   SIGNAL BU12543_D : STD_LOGIC;
   SIGNAL BU12543_CE : STD_LOGIC;
   SIGNAL BU12543_CLK : STD_LOGIC;
   SIGNAL BU12543_A0 : STD_LOGIC;
   SIGNAL BU12543_A1 : STD_LOGIC;
   SIGNAL BU12543_A2 : STD_LOGIC;
   SIGNAL BU12543_A3 : STD_LOGIC;
   SIGNAL BU12543_Q : STD_LOGIC;
   SIGNAL BU12544_D : STD_LOGIC;
   SIGNAL BU12544_CE : STD_LOGIC;
   SIGNAL BU12544_CLK : STD_LOGIC;
   SIGNAL BU12544_A0 : STD_LOGIC;
   SIGNAL BU12544_A1 : STD_LOGIC;
   SIGNAL BU12544_A2 : STD_LOGIC;
   SIGNAL BU12544_A3 : STD_LOGIC;
   SIGNAL BU12544_Q : STD_LOGIC;
   SIGNAL BU12545_D : STD_LOGIC;
   SIGNAL BU12545_CE : STD_LOGIC;
   SIGNAL BU12545_CLK : STD_LOGIC;
   SIGNAL BU12545_A0 : STD_LOGIC;
   SIGNAL BU12545_A1 : STD_LOGIC;
   SIGNAL BU12545_A2 : STD_LOGIC;
   SIGNAL BU12545_A3 : STD_LOGIC;
   SIGNAL BU12545_Q : STD_LOGIC;
   SIGNAL BU12546_D : STD_LOGIC;
   SIGNAL BU12546_CE : STD_LOGIC;
   SIGNAL BU12546_CLK : STD_LOGIC;
   SIGNAL BU12546_A0 : STD_LOGIC;
   SIGNAL BU12546_A1 : STD_LOGIC;
   SIGNAL BU12546_A2 : STD_LOGIC;
   SIGNAL BU12546_A3 : STD_LOGIC;
   SIGNAL BU12546_Q : STD_LOGIC;
   SIGNAL BU12547_D : STD_LOGIC;
   SIGNAL BU12547_CE : STD_LOGIC;
   SIGNAL BU12547_CLK : STD_LOGIC;
   SIGNAL BU12547_A0 : STD_LOGIC;
   SIGNAL BU12547_A1 : STD_LOGIC;
   SIGNAL BU12547_A2 : STD_LOGIC;
   SIGNAL BU12547_A3 : STD_LOGIC;
   SIGNAL BU12547_Q : STD_LOGIC;
   SIGNAL BU12548_D : STD_LOGIC;
   SIGNAL BU12548_CE : STD_LOGIC;
   SIGNAL BU12548_CLK : STD_LOGIC;
   SIGNAL BU12548_A0 : STD_LOGIC;
   SIGNAL BU12548_A1 : STD_LOGIC;
   SIGNAL BU12548_A2 : STD_LOGIC;
   SIGNAL BU12548_A3 : STD_LOGIC;
   SIGNAL BU12548_Q : STD_LOGIC;
   SIGNAL BU12549_D : STD_LOGIC;
   SIGNAL BU12549_CE : STD_LOGIC;
   SIGNAL BU12549_CLK : STD_LOGIC;
   SIGNAL BU12549_A0 : STD_LOGIC;
   SIGNAL BU12549_A1 : STD_LOGIC;
   SIGNAL BU12549_A2 : STD_LOGIC;
   SIGNAL BU12549_A3 : STD_LOGIC;
   SIGNAL BU12549_Q : STD_LOGIC;
   SIGNAL BU12550_Q : STD_LOGIC_VECTOR(3 DOWNTO 0);
   SIGNAL BU12550_CLK : STD_LOGIC;
   SIGNAL BU12550_UP : STD_LOGIC;
   SIGNAL BU12550_CE : STD_LOGIC;
   SIGNAL BU12579_I0 : STD_LOGIC;
   SIGNAL BU12579_I1 : STD_LOGIC;
   SIGNAL BU12579_I2 : STD_LOGIC;
   SIGNAL BU12579_I3 : STD_LOGIC;
   SIGNAL BU12579_O : STD_LOGIC;
   SIGNAL BU12583_I0 : STD_LOGIC;
   SIGNAL BU12583_I1 : STD_LOGIC;
   SIGNAL BU12583_I2 : STD_LOGIC;
   SIGNAL BU12583_I3 : STD_LOGIC;
   SIGNAL BU12583_O : STD_LOGIC;
   SIGNAL BU12584_D : STD_LOGIC;
   SIGNAL BU12584_C : STD_LOGIC;
   SIGNAL BU12584_CE : STD_LOGIC;
   SIGNAL BU12584_Q : STD_LOGIC;
   SIGNAL BU12587_I0 : STD_LOGIC;
   SIGNAL BU12587_I1 : STD_LOGIC;
   SIGNAL BU12587_I2 : STD_LOGIC;
   SIGNAL BU12587_I3 : STD_LOGIC;
   SIGNAL BU12587_O : STD_LOGIC;
   SIGNAL BU12588_ND : STD_LOGIC;
   SIGNAL BU12588_RDY : STD_LOGIC;
   SIGNAL BU12588_CLK : STD_LOGIC;
   SIGNAL BU12588_RFD : STD_LOGIC;
   SIGNAL BU12588_DIN : STD_LOGIC_VECTOR(25 DOWNTO 0);
   SIGNAL BU12588_DOUT : STD_LOGIC_VECTOR(42 DOWNTO 0);
   SIGNAL BU19118_I : STD_LOGIC_VECTOR(12 DOWNTO 0);
   SIGNAL BU19118_O : STD_LOGIC;
   SIGNAL BU19133_I0 : STD_LOGIC;
   SIGNAL BU19133_I1 : STD_LOGIC;
   SIGNAL BU19133_I2 : STD_LOGIC;
   SIGNAL BU19133_I3 : STD_LOGIC;
   SIGNAL BU19133_O : STD_LOGIC;
   SIGNAL BU19134_A : STD_LOGIC_VECTOR(29 DOWNTO 0);
   SIGNAL BU19134_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU19134_S : STD_LOGIC_VECTOR(30 DOWNTO 0);
   SIGNAL BU19259_I0 : STD_LOGIC;
   SIGNAL BU19259_I1 : STD_LOGIC;
   SIGNAL BU19259_I2 : STD_LOGIC;
   SIGNAL BU19259_I3 : STD_LOGIC;
   SIGNAL BU19259_O : STD_LOGIC;
   SIGNAL BU19261_I0 : STD_LOGIC;
   SIGNAL BU19261_I1 : STD_LOGIC;
   SIGNAL BU19261_I2 : STD_LOGIC;
   SIGNAL BU19261_I3 : STD_LOGIC;
   SIGNAL BU19261_O : STD_LOGIC;
   SIGNAL BU19262_D : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU19262_Q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU19262_CLK : STD_LOGIC;
   SIGNAL BU19262_SCLR : STD_LOGIC;
   SIGNAL BU19262_SSET : STD_LOGIC;
   SIGNAL BU19379_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU19379_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU19379_CLK : STD_LOGIC;
   SIGNAL BU19379_SCLR : STD_LOGIC;
   SIGNAL BU19379_SSET : STD_LOGIC;
   SIGNAL BU19386_D : STD_LOGIC;
   SIGNAL BU19386_C : STD_LOGIC;
   SIGNAL BU19386_CE : STD_LOGIC;
   SIGNAL BU19386_Q : STD_LOGIC;
   SIGNAL BU19389_ND : STD_LOGIC;
   SIGNAL BU19389_RDY : STD_LOGIC;
   SIGNAL BU19389_CLK : STD_LOGIC;
   SIGNAL BU19389_RFD : STD_LOGIC;
   SIGNAL BU19389_DIN : STD_LOGIC_VECTOR(29 DOWNTO 0);
   SIGNAL BU19389_SEL_O : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU19389_DOUT : STD_LOGIC_VECTOR(48 DOWNTO 0);
   SIGNAL BU25395_I0 : STD_LOGIC;
   SIGNAL BU25395_I1 : STD_LOGIC;
   SIGNAL BU25395_I2 : STD_LOGIC;
   SIGNAL BU25395_I3 : STD_LOGIC;
   SIGNAL BU25395_O : STD_LOGIC;
   SIGNAL BU25397_I0 : STD_LOGIC;
   SIGNAL BU25397_I1 : STD_LOGIC;
   SIGNAL BU25397_I2 : STD_LOGIC;
   SIGNAL BU25397_I3 : STD_LOGIC;
   SIGNAL BU25397_O : STD_LOGIC;
   SIGNAL BU25400_D : STD_LOGIC;
   SIGNAL BU25400_C : STD_LOGIC;
   SIGNAL BU25400_CE : STD_LOGIC;
   SIGNAL BU25400_Q : STD_LOGIC;
   SIGNAL BU25405_I : STD_LOGIC_VECTOR(18 DOWNTO 0);
   SIGNAL BU25405_O : STD_LOGIC;
   SIGNAL BU25427_I0 : STD_LOGIC;
   SIGNAL BU25427_I1 : STD_LOGIC;
   SIGNAL BU25427_I2 : STD_LOGIC;
   SIGNAL BU25427_I3 : STD_LOGIC;
   SIGNAL BU25427_O : STD_LOGIC;
   SIGNAL BU25428_A : STD_LOGIC_VECTOR(29 DOWNTO 0);
   SIGNAL BU25428_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU25428_S : STD_LOGIC_VECTOR(30 DOWNTO 0);
   SIGNAL BU25553_I0 : STD_LOGIC;
   SIGNAL BU25553_I1 : STD_LOGIC;
   SIGNAL BU25553_I2 : STD_LOGIC;
   SIGNAL BU25553_I3 : STD_LOGIC;
   SIGNAL BU25553_O : STD_LOGIC;
   SIGNAL BU25555_I0 : STD_LOGIC;
   SIGNAL BU25555_I1 : STD_LOGIC;
   SIGNAL BU25555_I2 : STD_LOGIC;
   SIGNAL BU25555_I3 : STD_LOGIC;
   SIGNAL BU25555_O : STD_LOGIC;
   SIGNAL BU25556_D : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU25556_Q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU25556_CLK : STD_LOGIC;
   SIGNAL BU25556_CE : STD_LOGIC;
   SIGNAL BU25556_SCLR : STD_LOGIC;
   SIGNAL BU25556_SSET : STD_LOGIC;
   SIGNAL BU25676_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU25676_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU25676_CLK : STD_LOGIC;
   SIGNAL BU25676_CE : STD_LOGIC;
   SIGNAL BU25676_SCLR : STD_LOGIC;
   SIGNAL BU25676_SSET : STD_LOGIC;
   SIGNAL BU25688_I : STD_LOGIC_VECTOR(18 DOWNTO 0);
   SIGNAL BU25688_O : STD_LOGIC;
   SIGNAL BU25710_I0 : STD_LOGIC;
   SIGNAL BU25710_I1 : STD_LOGIC;
   SIGNAL BU25710_I2 : STD_LOGIC;
   SIGNAL BU25710_I3 : STD_LOGIC;
   SIGNAL BU25710_O : STD_LOGIC;
   SIGNAL BU25711_A : STD_LOGIC_VECTOR(29 DOWNTO 0);
   SIGNAL BU25711_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU25711_S : STD_LOGIC_VECTOR(30 DOWNTO 0);
   SIGNAL BU25836_I0 : STD_LOGIC;
   SIGNAL BU25836_I1 : STD_LOGIC;
   SIGNAL BU25836_I2 : STD_LOGIC;
   SIGNAL BU25836_I3 : STD_LOGIC;
   SIGNAL BU25836_O : STD_LOGIC;
   SIGNAL BU25838_I0 : STD_LOGIC;
   SIGNAL BU25838_I1 : STD_LOGIC;
   SIGNAL BU25838_I2 : STD_LOGIC;
   SIGNAL BU25838_I3 : STD_LOGIC;
   SIGNAL BU25838_O : STD_LOGIC;
   SIGNAL BU25839_D : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU25839_Q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU25839_CLK : STD_LOGIC;
   SIGNAL BU25839_CE : STD_LOGIC;
   SIGNAL BU25839_SCLR : STD_LOGIC;
   SIGNAL BU25839_SSET : STD_LOGIC;
   SIGNAL BU25959_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU25959_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU25959_CLK : STD_LOGIC;
   SIGNAL BU25959_CE : STD_LOGIC;
   SIGNAL BU25959_SCLR : STD_LOGIC;
   SIGNAL BU25959_SSET : STD_LOGIC;
   SIGNAL n0 : STD_LOGIC := '0';
   SIGNAL n1 : STD_LOGIC := '1';
   SIGNAL n2 : STD_LOGIC;
   SIGNAL n3 : STD_LOGIC;
   SIGNAL n4 : STD_LOGIC;
   SIGNAL n5 : STD_LOGIC;
   SIGNAL n6 : STD_LOGIC;
   SIGNAL n7 : STD_LOGIC;
   SIGNAL n8 : STD_LOGIC;
   SIGNAL n9 : STD_LOGIC;
   SIGNAL n10 : STD_LOGIC;
   SIGNAL n11 : STD_LOGIC;
   SIGNAL n12 : STD_LOGIC;
   SIGNAL n13 : STD_LOGIC;
   SIGNAL n14 : STD_LOGIC;
   SIGNAL n15 : STD_LOGIC;
   SIGNAL n16 : STD_LOGIC;
   SIGNAL n17 : STD_LOGIC;
   SIGNAL n18 : STD_LOGIC;
   SIGNAL n19 : STD_LOGIC;
   SIGNAL n20 : STD_LOGIC;
   SIGNAL n21 : STD_LOGIC;
   SIGNAL n22 : STD_LOGIC;
   SIGNAL n23 : STD_LOGIC;
   SIGNAL n24 : STD_LOGIC;
   SIGNAL n25 : STD_LOGIC;
   SIGNAL n26 : STD_LOGIC;
   SIGNAL n27 : STD_LOGIC;
   SIGNAL n28 : STD_LOGIC;
   SIGNAL n29 : STD_LOGIC;
   SIGNAL n30 : STD_LOGIC;
   SIGNAL n31 : STD_LOGIC;
   SIGNAL n32 : STD_LOGIC;
   SIGNAL n33 : STD_LOGIC;
   SIGNAL n34 : STD_LOGIC;
   SIGNAL n35 : STD_LOGIC;
   SIGNAL n36 : STD_LOGIC;
   SIGNAL n37 : STD_LOGIC;
   SIGNAL n38 : STD_LOGIC;
   SIGNAL n39 : STD_LOGIC;
   SIGNAL n40 : STD_LOGIC;
   SIGNAL n41 : STD_LOGIC;
   SIGNAL n42 : STD_LOGIC;
   SIGNAL n43 : STD_LOGIC;
   SIGNAL n44 : STD_LOGIC;
   SIGNAL n45 : STD_LOGIC;
   SIGNAL n46 : STD_LOGIC;
   SIGNAL n47 : STD_LOGIC;
   SIGNAL n48 : STD_LOGIC;
   SIGNAL n49 : STD_LOGIC;
   SIGNAL n50 : STD_LOGIC;
   SIGNAL n54 : STD_LOGIC;
   SIGNAL n55 : STD_LOGIC;
   SIGNAL n58 : STD_LOGIC;
   SIGNAL n59 : STD_LOGIC;
   SIGNAL n60 : STD_LOGIC;
   SIGNAL n61 : STD_LOGIC;
   SIGNAL n62 : STD_LOGIC;
   SIGNAL n63 : STD_LOGIC;
   SIGNAL n64 : STD_LOGIC;
   SIGNAL n65 : STD_LOGIC;
   SIGNAL n66 : STD_LOGIC;
   SIGNAL n67 : STD_LOGIC;
   SIGNAL n68 : STD_LOGIC;
   SIGNAL n69 : STD_LOGIC;
   SIGNAL n70 : STD_LOGIC;
   SIGNAL n71 : STD_LOGIC;
   SIGNAL n72 : STD_LOGIC;
   SIGNAL n73 : STD_LOGIC;
   SIGNAL n74 : STD_LOGIC;
   SIGNAL n75 : STD_LOGIC;
   SIGNAL n76 : STD_LOGIC;
   SIGNAL n77 : STD_LOGIC;
   SIGNAL n78 : STD_LOGIC;
   SIGNAL n79 : STD_LOGIC;
   SIGNAL n80 : STD_LOGIC;
   SIGNAL n81 : STD_LOGIC;
   SIGNAL n82 : STD_LOGIC;
   SIGNAL n83 : STD_LOGIC;
   SIGNAL n84 : STD_LOGIC;
   SIGNAL n85 : STD_LOGIC;
   SIGNAL n86 : STD_LOGIC;
   SIGNAL n87 : STD_LOGIC;
   SIGNAL n88 : STD_LOGIC;
   SIGNAL n89 : STD_LOGIC;
   SIGNAL n90 : STD_LOGIC;
   SIGNAL n91 : STD_LOGIC;
   SIGNAL n92 : STD_LOGIC;
   SIGNAL n93 : STD_LOGIC;
   SIGNAL n94 : STD_LOGIC;
   SIGNAL n95 : STD_LOGIC;
   SIGNAL n96 : STD_LOGIC;
   SIGNAL n97 : STD_LOGIC;
   SIGNAL n98 : STD_LOGIC;
   SIGNAL n99 : STD_LOGIC;
   SIGNAL n100 : STD_LOGIC;
   SIGNAL n101 : STD_LOGIC;
   SIGNAL n102 : STD_LOGIC;
   SIGNAL n103 : STD_LOGIC;
   SIGNAL n104 : STD_LOGIC;
   SIGNAL n105 : STD_LOGIC;
   SIGNAL n106 : STD_LOGIC;
   SIGNAL n107 : STD_LOGIC;
   SIGNAL n108 : STD_LOGIC;
   SIGNAL n109 : STD_LOGIC;
   SIGNAL n110 : STD_LOGIC;
   SIGNAL n111 : STD_LOGIC;
   SIGNAL n112 : STD_LOGIC;
   SIGNAL n113 : STD_LOGIC;
   SIGNAL n114 : STD_LOGIC;
   SIGNAL n115 : STD_LOGIC;
   SIGNAL n116 : STD_LOGIC;
   SIGNAL n117 : STD_LOGIC;
   SIGNAL n118 : STD_LOGIC;
   SIGNAL n119 : STD_LOGIC;
   SIGNAL n120 : STD_LOGIC;
   SIGNAL n121 : STD_LOGIC;
   SIGNAL n122 : STD_LOGIC;
   SIGNAL n123 : STD_LOGIC;
   SIGNAL n124 : STD_LOGIC;
   SIGNAL n125 : STD_LOGIC;
   SIGNAL n126 : STD_LOGIC;
   SIGNAL n127 : STD_LOGIC;
   SIGNAL n128 : STD_LOGIC;
   SIGNAL n129 : STD_LOGIC;
   SIGNAL n130 : STD_LOGIC;
   SIGNAL n131 : STD_LOGIC;
   SIGNAL n132 : STD_LOGIC;
   SIGNAL n133 : STD_LOGIC;
   SIGNAL n134 : STD_LOGIC;
   SIGNAL n135 : STD_LOGIC;
   SIGNAL n136 : STD_LOGIC;
   SIGNAL n137 : STD_LOGIC;
   SIGNAL n138 : STD_LOGIC;
   SIGNAL n139 : STD_LOGIC;
   SIGNAL n140 : STD_LOGIC;
   SIGNAL n141 : STD_LOGIC;
   SIGNAL n142 : STD_LOGIC;
   SIGNAL n143 : STD_LOGIC;
   SIGNAL n144 : STD_LOGIC;
   SIGNAL n145 : STD_LOGIC;
   SIGNAL n146 : STD_LOGIC;
   SIGNAL n147 : STD_LOGIC;
   SIGNAL n148 : STD_LOGIC;
   SIGNAL n149 : STD_LOGIC;
   SIGNAL n150 : STD_LOGIC;
   SIGNAL n151 : STD_LOGIC;
   SIGNAL n152 : STD_LOGIC;
   SIGNAL n153 : STD_LOGIC;
   SIGNAL n154 : STD_LOGIC;
   SIGNAL n155 : STD_LOGIC;
   SIGNAL n156 : STD_LOGIC;
   SIGNAL n157 : STD_LOGIC;
   SIGNAL n158 : STD_LOGIC;
   SIGNAL n159 : STD_LOGIC;
   SIGNAL n160 : STD_LOGIC;
   SIGNAL n161 : STD_LOGIC;
   SIGNAL n162 : STD_LOGIC;
   SIGNAL n163 : STD_LOGIC;
   SIGNAL n164 : STD_LOGIC;
   SIGNAL n165 : STD_LOGIC;
   SIGNAL n166 : STD_LOGIC;
   SIGNAL n167 : STD_LOGIC;
   SIGNAL n168 : STD_LOGIC;
   SIGNAL n169 : STD_LOGIC;
   SIGNAL n170 : STD_LOGIC;
   SIGNAL n171 : STD_LOGIC;
   SIGNAL n172 : STD_LOGIC;
   SIGNAL n173 : STD_LOGIC;
   SIGNAL n174 : STD_LOGIC;
   SIGNAL n175 : STD_LOGIC;
   SIGNAL n176 : STD_LOGIC;
   SIGNAL n177 : STD_LOGIC;
   SIGNAL n178 : STD_LOGIC;
   SIGNAL n179 : STD_LOGIC;
   SIGNAL n180 : STD_LOGIC;
   SIGNAL n181 : STD_LOGIC;
   SIGNAL n182 : STD_LOGIC;
   SIGNAL n183 : STD_LOGIC;
   SIGNAL n184 : STD_LOGIC;
   SIGNAL n185 : STD_LOGIC;
   SIGNAL n186 : STD_LOGIC;
   SIGNAL n187 : STD_LOGIC;
   SIGNAL n188 : STD_LOGIC;
   SIGNAL n189 : STD_LOGIC;
   SIGNAL n190 : STD_LOGIC;
   SIGNAL n191 : STD_LOGIC;
   SIGNAL n192 : STD_LOGIC;
   SIGNAL n193 : STD_LOGIC;
   SIGNAL n194 : STD_LOGIC;
   SIGNAL n195 : STD_LOGIC;
   SIGNAL n196 : STD_LOGIC;
   SIGNAL n197 : STD_LOGIC;
   SIGNAL n198 : STD_LOGIC;
   SIGNAL n199 : STD_LOGIC;
   SIGNAL n200 : STD_LOGIC;
   SIGNAL n201 : STD_LOGIC;
   SIGNAL n202 : STD_LOGIC;
   SIGNAL n203 : STD_LOGIC;
   SIGNAL n204 : STD_LOGIC;
   SIGNAL n205 : STD_LOGIC;
   SIGNAL n206 : STD_LOGIC;
   SIGNAL n207 : STD_LOGIC;
   SIGNAL n208 : STD_LOGIC;
   SIGNAL n209 : STD_LOGIC;
   SIGNAL n210 : STD_LOGIC;
   SIGNAL n211 : STD_LOGIC;
   SIGNAL n212 : STD_LOGIC;
   SIGNAL n213 : STD_LOGIC;
   SIGNAL n214 : STD_LOGIC;
   SIGNAL n215 : STD_LOGIC;
   SIGNAL n216 : STD_LOGIC;
   SIGNAL n217 : STD_LOGIC;
   SIGNAL n218 : STD_LOGIC;
   SIGNAL n219 : STD_LOGIC;
   SIGNAL n220 : STD_LOGIC;
   SIGNAL n221 : STD_LOGIC;
   SIGNAL n222 : STD_LOGIC;
   SIGNAL n223 : STD_LOGIC;
   SIGNAL n224 : STD_LOGIC;
   SIGNAL n225 : STD_LOGIC;
   SIGNAL n226 : STD_LOGIC;
   SIGNAL n227 : STD_LOGIC;
   SIGNAL n228 : STD_LOGIC;
   SIGNAL n229 : STD_LOGIC;
   SIGNAL n230 : STD_LOGIC;
   SIGNAL n231 : STD_LOGIC;
   SIGNAL n232 : STD_LOGIC;
   SIGNAL n233 : STD_LOGIC;
   SIGNAL n234 : STD_LOGIC;
   SIGNAL n235 : STD_LOGIC;
   SIGNAL n236 : STD_LOGIC;
   SIGNAL n237 : STD_LOGIC;
   SIGNAL n238 : STD_LOGIC;
   SIGNAL n239 : STD_LOGIC;
   SIGNAL n240 : STD_LOGIC;
   SIGNAL n241 : STD_LOGIC;
   SIGNAL n242 : STD_LOGIC;
   SIGNAL n243 : STD_LOGIC;
   SIGNAL n244 : STD_LOGIC;
   SIGNAL n245 : STD_LOGIC;
   SIGNAL n246 : STD_LOGIC;
   SIGNAL n247 : STD_LOGIC;
   SIGNAL n248 : STD_LOGIC;
   SIGNAL n249 : STD_LOGIC;
   SIGNAL n250 : STD_LOGIC;
   SIGNAL n251 : STD_LOGIC;
   SIGNAL n252 : STD_LOGIC;
   SIGNAL n253 : STD_LOGIC;
   SIGNAL n254 : STD_LOGIC;
   SIGNAL n255 : STD_LOGIC;
   SIGNAL n256 : STD_LOGIC;
   SIGNAL n257 : STD_LOGIC;
   SIGNAL n258 : STD_LOGIC;
   SIGNAL n259 : STD_LOGIC;
   SIGNAL n260 : STD_LOGIC;
   SIGNAL n261 : STD_LOGIC;
   SIGNAL n262 : STD_LOGIC;
   SIGNAL n263 : STD_LOGIC;
   SIGNAL n264 : STD_LOGIC;
   SIGNAL n265 : STD_LOGIC;
   SIGNAL n266 : STD_LOGIC;
   SIGNAL n267 : STD_LOGIC;
   SIGNAL n268 : STD_LOGIC;
   SIGNAL n269 : STD_LOGIC;
   SIGNAL n270 : STD_LOGIC;
   SIGNAL n271 : STD_LOGIC;
   SIGNAL n272 : STD_LOGIC;
   SIGNAL n273 : STD_LOGIC;
   SIGNAL n274 : STD_LOGIC;
   SIGNAL n275 : STD_LOGIC;
   SIGNAL n276 : STD_LOGIC;
   SIGNAL n277 : STD_LOGIC;
   SIGNAL n278 : STD_LOGIC;
   SIGNAL n279 : STD_LOGIC;
   SIGNAL n280 : STD_LOGIC;
   SIGNAL n281 : STD_LOGIC;
   SIGNAL n282 : STD_LOGIC;
   SIGNAL n322 : STD_LOGIC;
   SIGNAL n369 : STD_LOGIC;
   SIGNAL n370 : STD_LOGIC;
   SIGNAL n371 : STD_LOGIC;
   SIGNAL n443 : STD_LOGIC;
   SIGNAL n444 : STD_LOGIC;
   SIGNAL n445 : STD_LOGIC;
   SIGNAL n446 : STD_LOGIC;
   SIGNAL n447 : STD_LOGIC;
   SIGNAL n448 : STD_LOGIC;
   SIGNAL n449 : STD_LOGIC;
   SIGNAL n450 : STD_LOGIC;
   SIGNAL n451 : STD_LOGIC;
   SIGNAL n452 : STD_LOGIC;
   SIGNAL n453 : STD_LOGIC;
   SIGNAL n454 : STD_LOGIC;
   SIGNAL n455 : STD_LOGIC;
   SIGNAL n456 : STD_LOGIC;
   SIGNAL n457 : STD_LOGIC;
   SIGNAL n488 : STD_LOGIC;
   SIGNAL n489 : STD_LOGIC;
   SIGNAL n490 : STD_LOGIC;
   SIGNAL n491 : STD_LOGIC;
   SIGNAL n492 : STD_LOGIC;
   SIGNAL n493 : STD_LOGIC;
   SIGNAL n494 : STD_LOGIC;
   SIGNAL n495 : STD_LOGIC;
   SIGNAL n496 : STD_LOGIC;
   SIGNAL n497 : STD_LOGIC;
   SIGNAL n498 : STD_LOGIC;
   SIGNAL n499 : STD_LOGIC;
   SIGNAL n500 : STD_LOGIC;
   SIGNAL n501 : STD_LOGIC;
   SIGNAL n502 : STD_LOGIC;
   SIGNAL n503 : STD_LOGIC;
   SIGNAL n504 : STD_LOGIC;
   SIGNAL n505 : STD_LOGIC;
   SIGNAL n506 : STD_LOGIC;
   SIGNAL n507 : STD_LOGIC;
   SIGNAL n508 : STD_LOGIC;
   SIGNAL n509 : STD_LOGIC;
   SIGNAL n510 : STD_LOGIC;
   SIGNAL n511 : STD_LOGIC;
   SIGNAL n512 : STD_LOGIC;
   SIGNAL n513 : STD_LOGIC;
   SIGNAL n514 : STD_LOGIC;
   SIGNAL n515 : STD_LOGIC;
   SIGNAL n516 : STD_LOGIC;
   SIGNAL n575 : STD_LOGIC;
   SIGNAL n605 : STD_LOGIC;
   SIGNAL n606 : STD_LOGIC;
   SIGNAL n607 : STD_LOGIC;
   SIGNAL n608 : STD_LOGIC;
   SIGNAL n609 : STD_LOGIC;
   SIGNAL n610 : STD_LOGIC;
   SIGNAL n611 : STD_LOGIC;
   SIGNAL n612 : STD_LOGIC;
   SIGNAL n613 : STD_LOGIC;
   SIGNAL n614 : STD_LOGIC;
   SIGNAL n615 : STD_LOGIC;
   SIGNAL n616 : STD_LOGIC;
   SIGNAL n617 : STD_LOGIC;
   SIGNAL n618 : STD_LOGIC;
   SIGNAL n647 : STD_LOGIC;
   SIGNAL n648 : STD_LOGIC;
   SIGNAL n649 : STD_LOGIC;
   SIGNAL n650 : STD_LOGIC;
   SIGNAL n651 : STD_LOGIC;
   SIGNAL n652 : STD_LOGIC;
   SIGNAL n653 : STD_LOGIC;
   SIGNAL n654 : STD_LOGIC;
   SIGNAL n655 : STD_LOGIC;
   SIGNAL n656 : STD_LOGIC;
   SIGNAL n657 : STD_LOGIC;
   SIGNAL n658 : STD_LOGIC;
   SIGNAL n659 : STD_LOGIC;
   SIGNAL n660 : STD_LOGIC;
   SIGNAL n661 : STD_LOGIC;
   SIGNAL n692 : STD_LOGIC;
   SIGNAL n693 : STD_LOGIC;
   SIGNAL n694 : STD_LOGIC;
   SIGNAL n695 : STD_LOGIC;
   SIGNAL n696 : STD_LOGIC;
   SIGNAL n697 : STD_LOGIC;
   SIGNAL n698 : STD_LOGIC;
   SIGNAL n699 : STD_LOGIC;
   SIGNAL n700 : STD_LOGIC;
   SIGNAL n701 : STD_LOGIC;
   SIGNAL n702 : STD_LOGIC;
   SIGNAL n703 : STD_LOGIC;
   SIGNAL n704 : STD_LOGIC;
   SIGNAL n705 : STD_LOGIC;
   SIGNAL n706 : STD_LOGIC;
   SIGNAL n707 : STD_LOGIC;
   SIGNAL n708 : STD_LOGIC;
   SIGNAL n709 : STD_LOGIC;
   SIGNAL n710 : STD_LOGIC;
   SIGNAL n711 : STD_LOGIC;
   SIGNAL n712 : STD_LOGIC;
   SIGNAL n713 : STD_LOGIC;
   SIGNAL n714 : STD_LOGIC;
   SIGNAL n715 : STD_LOGIC;
   SIGNAL n716 : STD_LOGIC;
   SIGNAL n717 : STD_LOGIC;
   SIGNAL n718 : STD_LOGIC;
   SIGNAL n719 : STD_LOGIC;
   SIGNAL n720 : STD_LOGIC;
   SIGNAL n955 : STD_LOGIC;
   SIGNAL n956 : STD_LOGIC;
   SIGNAL n957 : STD_LOGIC;
   SIGNAL n958 : STD_LOGIC;
   SIGNAL n959 : STD_LOGIC;
   SIGNAL n960 : STD_LOGIC;
   SIGNAL n961 : STD_LOGIC;
   SIGNAL n962 : STD_LOGIC;
   SIGNAL n963 : STD_LOGIC;
   SIGNAL n964 : STD_LOGIC;
   SIGNAL n965 : STD_LOGIC;
   SIGNAL n966 : STD_LOGIC;
   SIGNAL n967 : STD_LOGIC;
   SIGNAL n968 : STD_LOGIC;
   SIGNAL n1547 : STD_LOGIC;
   SIGNAL n1548 : STD_LOGIC;
   SIGNAL n1549 : STD_LOGIC;
   SIGNAL n1550 : STD_LOGIC;
   SIGNAL n1551 : STD_LOGIC;
   SIGNAL n1552 : STD_LOGIC;
   SIGNAL n1553 : STD_LOGIC;
   SIGNAL n1554 : STD_LOGIC;
   SIGNAL n1555 : STD_LOGIC;
   SIGNAL n1556 : STD_LOGIC;
   SIGNAL n1557 : STD_LOGIC;
   SIGNAL n1558 : STD_LOGIC;
   SIGNAL n1559 : STD_LOGIC;
   SIGNAL n1560 : STD_LOGIC;
   SIGNAL n1561 : STD_LOGIC;
   SIGNAL n1562 : STD_LOGIC;
   SIGNAL n1563 : STD_LOGIC;
   SIGNAL n1564 : STD_LOGIC;
   SIGNAL n1565 : STD_LOGIC;
   SIGNAL n1566 : STD_LOGIC;
   SIGNAL n1567 : STD_LOGIC;
   SIGNAL n1568 : STD_LOGIC;
   SIGNAL n1569 : STD_LOGIC;
   SIGNAL n1570 : STD_LOGIC;
   SIGNAL n1572 : STD_LOGIC;
   SIGNAL n1575 : STD_LOGIC;
   SIGNAL n1581 : STD_LOGIC;
   SIGNAL n1583 : STD_LOGIC;
   SIGNAL n2190 : STD_LOGIC;
   SIGNAL n2191 : STD_LOGIC;
   SIGNAL n2192 : STD_LOGIC;
   SIGNAL n2193 : STD_LOGIC;
   SIGNAL n2194 : STD_LOGIC;
   SIGNAL n2195 : STD_LOGIC;
   SIGNAL n2196 : STD_LOGIC;
   SIGNAL n2197 : STD_LOGIC;
   SIGNAL n2198 : STD_LOGIC;
   SIGNAL n2199 : STD_LOGIC;
   SIGNAL n2200 : STD_LOGIC;
   SIGNAL n2201 : STD_LOGIC;
   SIGNAL n2202 : STD_LOGIC;
   SIGNAL n2203 : STD_LOGIC;
   SIGNAL n2204 : STD_LOGIC;
   SIGNAL n2205 : STD_LOGIC;
   SIGNAL n2206 : STD_LOGIC;
   SIGNAL n2207 : STD_LOGIC;
   SIGNAL n2208 : STD_LOGIC;
   SIGNAL n2209 : STD_LOGIC;
   SIGNAL n2210 : STD_LOGIC;
   SIGNAL n2211 : STD_LOGIC;
   SIGNAL n2212 : STD_LOGIC;
   SIGNAL n2213 : STD_LOGIC;
   SIGNAL n2215 : STD_LOGIC;
   SIGNAL n2218 : STD_LOGIC;
   SIGNAL n2224 : STD_LOGIC;
   SIGNAL n2226 : STD_LOGIC;
   SIGNAL n2633 : STD_LOGIC;
   SIGNAL n2634 : STD_LOGIC;
   SIGNAL n2635 : STD_LOGIC;
   SIGNAL n2636 : STD_LOGIC;
   SIGNAL n2637 : STD_LOGIC;
   SIGNAL n2638 : STD_LOGIC;
   SIGNAL n2639 : STD_LOGIC;
   SIGNAL n2640 : STD_LOGIC;
   SIGNAL n2641 : STD_LOGIC;
   SIGNAL n2642 : STD_LOGIC;
   SIGNAL n2643 : STD_LOGIC;
   SIGNAL n2644 : STD_LOGIC;
   SIGNAL n2645 : STD_LOGIC;
   SIGNAL n2646 : STD_LOGIC;
   SIGNAL n2647 : STD_LOGIC;
   SIGNAL n2648 : STD_LOGIC;
   SIGNAL n2649 : STD_LOGIC;
   SIGNAL n2650 : STD_LOGIC;
   SIGNAL n2651 : STD_LOGIC;
   SIGNAL n2652 : STD_LOGIC;
   SIGNAL n2653 : STD_LOGIC;
   SIGNAL n2654 : STD_LOGIC;
   SIGNAL n2655 : STD_LOGIC;
   SIGNAL n2656 : STD_LOGIC;
   SIGNAL n2657 : STD_LOGIC;
   SIGNAL n2658 : STD_LOGIC;
   SIGNAL n2659 : STD_LOGIC;
   SIGNAL n2660 : STD_LOGIC;
   SIGNAL n2661 : STD_LOGIC;
   SIGNAL n2662 : STD_LOGIC;
   SIGNAL n2663 : STD_LOGIC;
   SIGNAL n2664 : STD_LOGIC;
   SIGNAL n2665 : STD_LOGIC;
   SIGNAL n2666 : STD_LOGIC;
   SIGNAL n2667 : STD_LOGIC;
   SIGNAL n2668 : STD_LOGIC;
   SIGNAL n2669 : STD_LOGIC;
   SIGNAL n2670 : STD_LOGIC;
   SIGNAL n2671 : STD_LOGIC;
   SIGNAL n2672 : STD_LOGIC;
   SIGNAL n2673 : STD_LOGIC;
   SIGNAL n2674 : STD_LOGIC;
   SIGNAL n2675 : STD_LOGIC;
   SIGNAL n2676 : STD_LOGIC;
   SIGNAL n2677 : STD_LOGIC;
   SIGNAL n2678 : STD_LOGIC;
   SIGNAL n2679 : STD_LOGIC;
   SIGNAL n2680 : STD_LOGIC;
   SIGNAL n2681 : STD_LOGIC;
   SIGNAL n2682 : STD_LOGIC;
   SIGNAL n2683 : STD_LOGIC;
   SIGNAL n2684 : STD_LOGIC;
   SIGNAL n2685 : STD_LOGIC;
   SIGNAL n2686 : STD_LOGIC;
   SIGNAL n2687 : STD_LOGIC;
   SIGNAL n2688 : STD_LOGIC;
   SIGNAL n2689 : STD_LOGIC;
   SIGNAL n2690 : STD_LOGIC;
   SIGNAL n2691 : STD_LOGIC;
   SIGNAL n2692 : STD_LOGIC;
   SIGNAL n2693 : STD_LOGIC;
   SIGNAL n2694 : STD_LOGIC;
   SIGNAL n2695 : STD_LOGIC;
   SIGNAL n2696 : STD_LOGIC;
   SIGNAL n2697 : STD_LOGIC;
   SIGNAL n2698 : STD_LOGIC;
   SIGNAL n2699 : STD_LOGIC;
   SIGNAL n2700 : STD_LOGIC;
   SIGNAL n2701 : STD_LOGIC;
   SIGNAL n2702 : STD_LOGIC;
   SIGNAL n2703 : STD_LOGIC;
   SIGNAL n2704 : STD_LOGIC;
   SIGNAL n2705 : STD_LOGIC;
   SIGNAL n2706 : STD_LOGIC;
   SIGNAL n2707 : STD_LOGIC;
   SIGNAL n2708 : STD_LOGIC;
   SIGNAL n2709 : STD_LOGIC;
   SIGNAL n2710 : STD_LOGIC;
   SIGNAL n2711 : STD_LOGIC;
   SIGNAL n2712 : STD_LOGIC;
   SIGNAL n2713 : STD_LOGIC;
   SIGNAL n2714 : STD_LOGIC;
   SIGNAL n2715 : STD_LOGIC;
   SIGNAL n2716 : STD_LOGIC;
   SIGNAL n2717 : STD_LOGIC;
   SIGNAL n2718 : STD_LOGIC;
   SIGNAL n2719 : STD_LOGIC;
   SIGNAL n2720 : STD_LOGIC;
   SIGNAL n2721 : STD_LOGIC;
   SIGNAL n2722 : STD_LOGIC;
   SIGNAL n2723 : STD_LOGIC;
   SIGNAL n2724 : STD_LOGIC;
   SIGNAL n2725 : STD_LOGIC;
   SIGNAL n2726 : STD_LOGIC;
   SIGNAL n2727 : STD_LOGIC;
   SIGNAL n2728 : STD_LOGIC;
   SIGNAL n2729 : STD_LOGIC;
   SIGNAL n2730 : STD_LOGIC;
   SIGNAL n2731 : STD_LOGIC;
   SIGNAL n2732 : STD_LOGIC;
   SIGNAL n2733 : STD_LOGIC;
   SIGNAL n2734 : STD_LOGIC;
   SIGNAL n2735 : STD_LOGIC;
   SIGNAL n2736 : STD_LOGIC;
   SIGNAL n2737 : STD_LOGIC;
   SIGNAL n2738 : STD_LOGIC;
   SIGNAL n2739 : STD_LOGIC;
   SIGNAL n2740 : STD_LOGIC;
   SIGNAL n2741 : STD_LOGIC;
   SIGNAL n2742 : STD_LOGIC;
   SIGNAL n2743 : STD_LOGIC;
   SIGNAL n2744 : STD_LOGIC;
   SIGNAL n2745 : STD_LOGIC;
   SIGNAL n2746 : STD_LOGIC;
   SIGNAL n2747 : STD_LOGIC;
   SIGNAL n2748 : STD_LOGIC;
   SIGNAL n2749 : STD_LOGIC;
   SIGNAL n2750 : STD_LOGIC;
   SIGNAL n2751 : STD_LOGIC;
   SIGNAL n2752 : STD_LOGIC;
   SIGNAL n2753 : STD_LOGIC;
   SIGNAL n2754 : STD_LOGIC;
   SIGNAL n2755 : STD_LOGIC;
   SIGNAL n2756 : STD_LOGIC;
   SIGNAL n2757 : STD_LOGIC;
   SIGNAL n2758 : STD_LOGIC;
   SIGNAL n2759 : STD_LOGIC;
   SIGNAL n2760 : STD_LOGIC;
   SIGNAL n2761 : STD_LOGIC;
   SIGNAL n2762 : STD_LOGIC;
   SIGNAL n2763 : STD_LOGIC;
   SIGNAL n2764 : STD_LOGIC;
   SIGNAL n2765 : STD_LOGIC;
   SIGNAL n2766 : STD_LOGIC;
   SIGNAL n2767 : STD_LOGIC;
   SIGNAL n2768 : STD_LOGIC;
   SIGNAL n2769 : STD_LOGIC;
   SIGNAL n2770 : STD_LOGIC;
   SIGNAL n2771 : STD_LOGIC;
   SIGNAL n2772 : STD_LOGIC;
   SIGNAL n2773 : STD_LOGIC;
   SIGNAL n2774 : STD_LOGIC;
   SIGNAL n2775 : STD_LOGIC;
   SIGNAL n2776 : STD_LOGIC;
   SIGNAL n2777 : STD_LOGIC;
   SIGNAL n2778 : STD_LOGIC;
   SIGNAL n2779 : STD_LOGIC;
   SIGNAL n2780 : STD_LOGIC;
   SIGNAL n2781 : STD_LOGIC;
   SIGNAL n2782 : STD_LOGIC;
   SIGNAL n2783 : STD_LOGIC;
   SIGNAL n2784 : STD_LOGIC;
   SIGNAL n2785 : STD_LOGIC;
   SIGNAL n2786 : STD_LOGIC;
   SIGNAL n2787 : STD_LOGIC;
   SIGNAL n2788 : STD_LOGIC;
   SIGNAL n2789 : STD_LOGIC;
   SIGNAL n2790 : STD_LOGIC;
   SIGNAL n2791 : STD_LOGIC;
   SIGNAL n2792 : STD_LOGIC;
   SIGNAL n2793 : STD_LOGIC;
   SIGNAL n2794 : STD_LOGIC;
   SIGNAL n2795 : STD_LOGIC;
   SIGNAL n2796 : STD_LOGIC;
   SIGNAL n2797 : STD_LOGIC;
   SIGNAL n2798 : STD_LOGIC;
   SIGNAL n2799 : STD_LOGIC;
   SIGNAL n2800 : STD_LOGIC;
   SIGNAL n2801 : STD_LOGIC;
   SIGNAL n3042 : STD_LOGIC;
   SIGNAL n3043 : STD_LOGIC;
   SIGNAL n3044 : STD_LOGIC;
   SIGNAL n3045 : STD_LOGIC;
   SIGNAL n3046 : STD_LOGIC;
   SIGNAL n3047 : STD_LOGIC;
   SIGNAL n3048 : STD_LOGIC;
   SIGNAL n3049 : STD_LOGIC;
   SIGNAL n3050 : STD_LOGIC;
   SIGNAL n3051 : STD_LOGIC;
   SIGNAL n3052 : STD_LOGIC;
   SIGNAL n3053 : STD_LOGIC;
   SIGNAL n3054 : STD_LOGIC;
   SIGNAL n3055 : STD_LOGIC;
   SIGNAL n3056 : STD_LOGIC;
   SIGNAL n3057 : STD_LOGIC;
   SIGNAL n3058 : STD_LOGIC;
   SIGNAL n3059 : STD_LOGIC;
   SIGNAL n3060 : STD_LOGIC;
   SIGNAL n3061 : STD_LOGIC;
   SIGNAL n3062 : STD_LOGIC;
   SIGNAL n3063 : STD_LOGIC;
   SIGNAL n3064 : STD_LOGIC;
   SIGNAL n3065 : STD_LOGIC;
   SIGNAL n3067 : STD_LOGIC;
   SIGNAL n3070 : STD_LOGIC;
   SIGNAL n3094 : STD_LOGIC;
   SIGNAL n3096 : STD_LOGIC;
   SIGNAL n3559 : STD_LOGIC;
   SIGNAL n3560 : STD_LOGIC;
   SIGNAL n3561 : STD_LOGIC;
   SIGNAL n3562 : STD_LOGIC;
   SIGNAL n3563 : STD_LOGIC;
   SIGNAL n3564 : STD_LOGIC;
   SIGNAL n3565 : STD_LOGIC;
   SIGNAL n3566 : STD_LOGIC;
   SIGNAL n3567 : STD_LOGIC;
   SIGNAL n3568 : STD_LOGIC;
   SIGNAL n3569 : STD_LOGIC;
   SIGNAL n3570 : STD_LOGIC;
   SIGNAL n3571 : STD_LOGIC;
   SIGNAL n3572 : STD_LOGIC;
   SIGNAL n3573 : STD_LOGIC;
   SIGNAL n3574 : STD_LOGIC;
   SIGNAL n3575 : STD_LOGIC;
   SIGNAL n3576 : STD_LOGIC;
   SIGNAL n3577 : STD_LOGIC;
   SIGNAL n3578 : STD_LOGIC;
   SIGNAL n3579 : STD_LOGIC;
   SIGNAL n3580 : STD_LOGIC;
   SIGNAL n3581 : STD_LOGIC;
   SIGNAL n3582 : STD_LOGIC;
   SIGNAL n3584 : STD_LOGIC;
   SIGNAL n3587 : STD_LOGIC;
   SIGNAL n3611 : STD_LOGIC;
   SIGNAL n3613 : STD_LOGIC;
   SIGNAL n4473 : STD_LOGIC;
   SIGNAL n6719 : STD_LOGIC;
   SIGNAL n6720 : STD_LOGIC;
   SIGNAL n6721 : STD_LOGIC;
   SIGNAL n6722 : STD_LOGIC;
   SIGNAL n6723 : STD_LOGIC;
   SIGNAL n6724 : STD_LOGIC;
   SIGNAL n6725 : STD_LOGIC;
   SIGNAL n6726 : STD_LOGIC;
   SIGNAL n6727 : STD_LOGIC;
   SIGNAL n6728 : STD_LOGIC;
   SIGNAL n6729 : STD_LOGIC;
   SIGNAL n6730 : STD_LOGIC;
   SIGNAL n6731 : STD_LOGIC;
   SIGNAL n6732 : STD_LOGIC;
   SIGNAL n6733 : STD_LOGIC;
   SIGNAL n6734 : STD_LOGIC;
   SIGNAL n6735 : STD_LOGIC;
   SIGNAL n6736 : STD_LOGIC;
   SIGNAL n6737 : STD_LOGIC;
   SIGNAL n6738 : STD_LOGIC;
   SIGNAL n6739 : STD_LOGIC;
   SIGNAL n6740 : STD_LOGIC;
   SIGNAL n6741 : STD_LOGIC;
   SIGNAL n6742 : STD_LOGIC;
   SIGNAL n6743 : STD_LOGIC;
   SIGNAL n6744 : STD_LOGIC;
   SIGNAL n6745 : STD_LOGIC;
   SIGNAL n6746 : STD_LOGIC;
   SIGNAL n6747 : STD_LOGIC;
   SIGNAL n6748 : STD_LOGIC;
   SIGNAL n6749 : STD_LOGIC;
   SIGNAL n6750 : STD_LOGIC;
   SIGNAL n6751 : STD_LOGIC;
   SIGNAL n6752 : STD_LOGIC;
   SIGNAL n6753 : STD_LOGIC;
   SIGNAL n6754 : STD_LOGIC;
   SIGNAL n6755 : STD_LOGIC;
   SIGNAL n6756 : STD_LOGIC;
   SIGNAL n6757 : STD_LOGIC;
   SIGNAL n6758 : STD_LOGIC;
   SIGNAL n6759 : STD_LOGIC;
   SIGNAL n6760 : STD_LOGIC;
   SIGNAL n6761 : STD_LOGIC;
   SIGNAL n6762 : STD_LOGIC;
   SIGNAL n6763 : STD_LOGIC;
   SIGNAL n6764 : STD_LOGIC;
   SIGNAL n6765 : STD_LOGIC;
   SIGNAL n6766 : STD_LOGIC;
   SIGNAL n6767 : STD_LOGIC;
   SIGNAL n6768 : STD_LOGIC;
   SIGNAL n6769 : STD_LOGIC;
   SIGNAL n6770 : STD_LOGIC;
   SIGNAL n6771 : STD_LOGIC;
   SIGNAL n6772 : STD_LOGIC;
   SIGNAL n6773 : STD_LOGIC;
   SIGNAL n6774 : STD_LOGIC;
   SIGNAL n6775 : STD_LOGIC;
   SIGNAL n6776 : STD_LOGIC;
   SIGNAL n6777 : STD_LOGIC;
   SIGNAL n6778 : STD_LOGIC;
   SIGNAL n6779 : STD_LOGIC;
   SIGNAL n6780 : STD_LOGIC;
   SIGNAL n6781 : STD_LOGIC;
   SIGNAL n6782 : STD_LOGIC;
   SIGNAL n6783 : STD_LOGIC;
   SIGNAL n6784 : STD_LOGIC;
   SIGNAL n6785 : STD_LOGIC;
   SIGNAL n6786 : STD_LOGIC;
   SIGNAL n6787 : STD_LOGIC;
   SIGNAL n6788 : STD_LOGIC;
   SIGNAL n6789 : STD_LOGIC;
   SIGNAL n6790 : STD_LOGIC;
   SIGNAL n6791 : STD_LOGIC;
   SIGNAL n6857 : STD_LOGIC;
   SIGNAL n6858 : STD_LOGIC;
   SIGNAL n6859 : STD_LOGIC;
   SIGNAL n6860 : STD_LOGIC;
   SIGNAL n6861 : STD_LOGIC;
   SIGNAL n6862 : STD_LOGIC;
   SIGNAL n6863 : STD_LOGIC;
   SIGNAL n7206 : STD_LOGIC;
   SIGNAL n7333 : STD_LOGIC;
   SIGNAL n7334 : STD_LOGIC;
   SIGNAL n7335 : STD_LOGIC;
   SIGNAL n7336 : STD_LOGIC;
   SIGNAL n7337 : STD_LOGIC;
   SIGNAL n7338 : STD_LOGIC;
   SIGNAL n7339 : STD_LOGIC;
   SIGNAL n7340 : STD_LOGIC;
   SIGNAL n7341 : STD_LOGIC;
   SIGNAL n7342 : STD_LOGIC;
   SIGNAL n7343 : STD_LOGIC;
   SIGNAL n7344 : STD_LOGIC;
   SIGNAL n7345 : STD_LOGIC;
   SIGNAL n7346 : STD_LOGIC;
   SIGNAL n7347 : STD_LOGIC;
   SIGNAL n7348 : STD_LOGIC;
   SIGNAL n7349 : STD_LOGIC;
   SIGNAL n7350 : STD_LOGIC;
   SIGNAL n7351 : STD_LOGIC;
   SIGNAL n7352 : STD_LOGIC;
   SIGNAL n7353 : STD_LOGIC;
   SIGNAL n7354 : STD_LOGIC;
   SIGNAL n7355 : STD_LOGIC;
   SIGNAL n7356 : STD_LOGIC;
   SIGNAL n7357 : STD_LOGIC;
   SIGNAL n7358 : STD_LOGIC;
   SIGNAL n7359 : STD_LOGIC;
   SIGNAL n7360 : STD_LOGIC;
   SIGNAL n7361 : STD_LOGIC;
   SIGNAL n7362 : STD_LOGIC;
   SIGNAL n7364 : STD_LOGIC;
   SIGNAL n7367 : STD_LOGIC;
   SIGNAL n7381 : STD_LOGIC;
   SIGNAL n7383 : STD_LOGIC;
   SIGNAL n8099 : STD_LOGIC;
   SIGNAL n8100 : STD_LOGIC;
   SIGNAL n8101 : STD_LOGIC;
   SIGNAL n8102 : STD_LOGIC;
   SIGNAL n8103 : STD_LOGIC;
   SIGNAL n8104 : STD_LOGIC;
   SIGNAL n8105 : STD_LOGIC;
   SIGNAL n8106 : STD_LOGIC;
   SIGNAL n8107 : STD_LOGIC;
   SIGNAL n8108 : STD_LOGIC;
   SIGNAL n8109 : STD_LOGIC;
   SIGNAL n8110 : STD_LOGIC;
   SIGNAL n8111 : STD_LOGIC;
   SIGNAL n8112 : STD_LOGIC;
   SIGNAL n8113 : STD_LOGIC;
   SIGNAL n8114 : STD_LOGIC;
   SIGNAL n8115 : STD_LOGIC;
   SIGNAL n8116 : STD_LOGIC;
   SIGNAL n8117 : STD_LOGIC;
   SIGNAL n8118 : STD_LOGIC;
   SIGNAL n8119 : STD_LOGIC;
   SIGNAL n8120 : STD_LOGIC;
   SIGNAL n8121 : STD_LOGIC;
   SIGNAL n8122 : STD_LOGIC;
   SIGNAL n8123 : STD_LOGIC;
   SIGNAL n8124 : STD_LOGIC;
   SIGNAL n8125 : STD_LOGIC;
   SIGNAL n8126 : STD_LOGIC;
   SIGNAL n8127 : STD_LOGIC;
   SIGNAL n8128 : STD_LOGIC;
   SIGNAL n8130 : STD_LOGIC;
   SIGNAL n8133 : STD_LOGIC;
   SIGNAL n8153 : STD_LOGIC;
   SIGNAL n8155 : STD_LOGIC;
   SIGNAL n8701 : STD_LOGIC;
   SIGNAL n8702 : STD_LOGIC;
   SIGNAL n8703 : STD_LOGIC;
   SIGNAL n8704 : STD_LOGIC;
   SIGNAL n8705 : STD_LOGIC;
   SIGNAL n8706 : STD_LOGIC;
   SIGNAL n8707 : STD_LOGIC;
   SIGNAL n8708 : STD_LOGIC;
   SIGNAL n8709 : STD_LOGIC;
   SIGNAL n8710 : STD_LOGIC;
   SIGNAL n8711 : STD_LOGIC;
   SIGNAL n8712 : STD_LOGIC;
   SIGNAL n8713 : STD_LOGIC;
   SIGNAL n8714 : STD_LOGIC;
   SIGNAL n8715 : STD_LOGIC;
   SIGNAL n8716 : STD_LOGIC;
   SIGNAL n8717 : STD_LOGIC;
   SIGNAL n8718 : STD_LOGIC;
   SIGNAL n8719 : STD_LOGIC;
   SIGNAL n8720 : STD_LOGIC;
   SIGNAL n8721 : STD_LOGIC;
   SIGNAL n8722 : STD_LOGIC;
   SIGNAL n8723 : STD_LOGIC;
   SIGNAL n8724 : STD_LOGIC;
   SIGNAL n8725 : STD_LOGIC;
   SIGNAL n8726 : STD_LOGIC;
   SIGNAL n8727 : STD_LOGIC;
   SIGNAL n8728 : STD_LOGIC;
   SIGNAL n8729 : STD_LOGIC;
   SIGNAL n8730 : STD_LOGIC;
   SIGNAL n8732 : STD_LOGIC;
   SIGNAL n8735 : STD_LOGIC;
   SIGNAL n8755 : STD_LOGIC;
   SIGNAL n8757 : STD_LOGIC;

BEGIN

   n166 <= DIN(0);
   n167 <= DIN(1);
   n168 <= DIN(2);
   n169 <= DIN(3);
   n170 <= DIN(4);
   n171 <= DIN(5);
   n172 <= DIN(6);
   n173 <= DIN(7);
   n174 <= DIN(8);
   n175 <= DIN(9);
   n176 <= DIN(10);
   n177 <= DIN(11);
   n178 <= DIN(12);
   n179 <= DIN(13);
   n180 <= ND;
   n183 <= CLK;
   n184 <= ADDR(0);
   n185 <= ADDR(1);
   n186 <= ADDR(2);
   n187 <= ADDR(3);
   n188 <= ADDR(4);
   n189 <= LD_DIN(0);
   n190 <= LD_DIN(1);
   n191 <= LD_DIN(2);
   n192 <= LD_DIN(3);
   n193 <= LD_DIN(4);
   n194 <= LD_DIN(5);
   n195 <= LD_DIN(6);
   n196 <= LD_DIN(7);
   n197 <= LD_DIN(8);
   n198 <= LD_DIN(9);
   n199 <= LD_DIN(10);
   n200 <= LD_DIN(11);
   n201 <= LD_DIN(12);
   n202 <= LD_DIN(13);
   n203 <= LD_DIN(14);
   n204 <= LD_DIN(15);
   n205 <= LD_DIN(16);
   n206 <= LD_DIN(17);
   n207 <= LD_DIN(18);
   n208 <= LD_DIN(19);
   n209 <= LD_DIN(20);
   n210 <= LD_DIN(21);
   n211 <= LD_DIN(22);
   n212 <= LD_DIN(23);
   n213 <= LD_DIN(24);
   n214 <= LD_DIN(25);
   n215 <= LD_DIN(26);
   n216 <= LD_DIN(27);
   n217 <= LD_DIN(28);
   n218 <= LD_DIN(29);
   n219 <= LD_DIN(30);
   n220 <= LD_DIN(31);
   n221 <= WE;
   n222 <= SEL;
   RDY <= n181;
   RFD <= n182;
   DOUT_I(0) <= n223;
   DOUT_I(1) <= n224;
   DOUT_I(2) <= n225;
   DOUT_I(3) <= n226;
   DOUT_I(4) <= n227;
   DOUT_I(5) <= n228;
   DOUT_I(6) <= n229;
   DOUT_I(7) <= n230;
   DOUT_I(8) <= n231;
   DOUT_I(9) <= n232;
   DOUT_I(10) <= n233;
   DOUT_I(11) <= n234;
   DOUT_I(12) <= n235;
   DOUT_I(13) <= n236;
   DOUT_I(14) <= n237;
   DOUT_I(15) <= n238;
   DOUT_I(16) <= n239;
   DOUT_I(17) <= n240;
   DOUT_I(18) <= n241;
   DOUT_I(19) <= n242;
   DOUT_I(20) <= n243;
   DOUT_I(21) <= n244;
   DOUT_I(22) <= n245;
   DOUT_I(23) <= n246;
   DOUT_I(24) <= n247;
   DOUT_I(25) <= n248;
   DOUT_I(26) <= n249;
   DOUT_I(27) <= n250;
   DOUT_I(28) <= n251;
   DOUT_I(29) <= n252;
   DOUT_Q(0) <= n253;
   DOUT_Q(1) <= n254;
   DOUT_Q(2) <= n255;
   DOUT_Q(3) <= n256;
   DOUT_Q(4) <= n257;
   DOUT_Q(5) <= n258;
   DOUT_Q(6) <= n259;
   DOUT_Q(7) <= n260;
   DOUT_Q(8) <= n261;
   DOUT_Q(9) <= n262;
   DOUT_Q(10) <= n263;
   DOUT_Q(11) <= n264;
   DOUT_Q(12) <= n265;
   DOUT_Q(13) <= n266;
   DOUT_Q(14) <= n267;
   DOUT_Q(15) <= n268;
   DOUT_Q(16) <= n269;
   DOUT_Q(17) <= n270;
   DOUT_Q(18) <= n271;
   DOUT_Q(19) <= n272;
   DOUT_Q(20) <= n273;
   DOUT_Q(21) <= n274;
   DOUT_Q(22) <= n275;
   DOUT_Q(23) <= n276;
   DOUT_Q(24) <= n277;
   DOUT_Q(25) <= n278;
   DOUT_Q(26) <= n279;
   DOUT_Q(27) <= n280;
   DOUT_Q(28) <= n281;
   DOUT_Q(29) <= n282;

   BU4_I0 <= n188;
   BU4_I1 <= n187;
   BU4_I2 <= n186;
   BU4_I3 <= n222;
   n54 <= BU4_O;
   BU4 : LUT4
      GENERIC MAP (
         INIT  => X"1000"
      )
      PORT MAP (
         I0 => BU4_I0,
         I1 => BU4_I1,
         I2 => BU4_I2,
         I3 => BU4_I3,
         O => BU4_O
      );

   BU8_I0 <= n54;
   BU8_I1 <= n221;
   BU8_I2 <= n185;
   BU8_I3 <= n184;
   n322 <= BU8_O;
   BU8 : LUT4
      GENERIC MAP (
         INIT  => X"0080"
      )
      PORT MAP (
         I0 => BU8_I0,
         I1 => BU8_I1,
         I2 => BU8_I2,
         I3 => BU8_I3,
         O => BU8_O
      );

   BU10_I0 <= '1';
   BU10_I1 <= '0';
   BU10_I2 <= '0';
   BU10_I3 <= '0';
   n182 <= BU10_O;
   BU10 : LUT4
      GENERIC MAP (
         INIT  => X"aaaa"
      )
      PORT MAP (
         I0 => BU10_I0,
         I1 => BU10_I1,
         I2 => BU10_I2,
         I3 => BU10_I3,
         O => BU10_O
      );

   BU1292_D <= n180;
   BU1292_C <= n183;
   BU1292_CE <= '1';
   n371 <= BU1292_Q;
   BU1292 : FDE
      PORT MAP (
         D => BU1292_D,
         C => BU1292_C,
         CE => BU1292_CE,
         Q => BU1292_Q
      );

   BU14_D <= n166;
   BU14_CE <= n180;
   BU14_CLK <= n183;
   BU14_A0 <= '0';
   BU14_A1 <= '1';
   BU14_A2 <= '0';
   BU14_A3 <= '0';
   n955 <= BU14_Q;
   BU14 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU14_D,
         CE => BU14_CE,
         CLK => BU14_CLK,
         A0 => BU14_A0,
         A1 => BU14_A1,
         A2 => BU14_A2,
         A3 => BU14_A3,
         Q => BU14_Q
      );

   BU16_D <= n955;
   BU16_C <= n183;
   BU16_CE <= n180;
   n618 <= BU16_Q;
   BU16 : FDE
      PORT MAP (
         D => BU16_D,
         C => BU16_C,
         CE => BU16_CE,
         Q => BU16_Q
      );

   BU17_D <= n167;
   BU17_CE <= n180;
   BU17_CLK <= n183;
   BU17_A0 <= '0';
   BU17_A1 <= '1';
   BU17_A2 <= '0';
   BU17_A3 <= '0';
   n956 <= BU17_Q;
   BU17 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU17_D,
         CE => BU17_CE,
         CLK => BU17_CLK,
         A0 => BU17_A0,
         A1 => BU17_A1,
         A2 => BU17_A2,
         A3 => BU17_A3,
         Q => BU17_Q
      );

   BU19_D <= n956;
   BU19_C <= n183;
   BU19_CE <= n180;
   n617 <= BU19_Q;
   BU19 : FDE
      PORT MAP (
         D => BU19_D,
         C => BU19_C,
         CE => BU19_CE,
         Q => BU19_Q
      );

   BU20_D <= n168;
   BU20_CE <= n180;
   BU20_CLK <= n183;
   BU20_A0 <= '0';
   BU20_A1 <= '1';
   BU20_A2 <= '0';
   BU20_A3 <= '0';
   n957 <= BU20_Q;
   BU20 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU20_D,
         CE => BU20_CE,
         CLK => BU20_CLK,
         A0 => BU20_A0,
         A1 => BU20_A1,
         A2 => BU20_A2,
         A3 => BU20_A3,
         Q => BU20_Q
      );

   BU22_D <= n957;
   BU22_C <= n183;
   BU22_CE <= n180;
   n616 <= BU22_Q;
   BU22 : FDE
      PORT MAP (
         D => BU22_D,
         C => BU22_C,
         CE => BU22_CE,
         Q => BU22_Q
      );

   BU23_D <= n169;
   BU23_CE <= n180;
   BU23_CLK <= n183;
   BU23_A0 <= '0';
   BU23_A1 <= '1';
   BU23_A2 <= '0';
   BU23_A3 <= '0';
   n958 <= BU23_Q;
   BU23 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU23_D,
         CE => BU23_CE,
         CLK => BU23_CLK,
         A0 => BU23_A0,
         A1 => BU23_A1,
         A2 => BU23_A2,
         A3 => BU23_A3,
         Q => BU23_Q
      );

   BU25_D <= n958;
   BU25_C <= n183;
   BU25_CE <= n180;
   n615 <= BU25_Q;
   BU25 : FDE
      PORT MAP (
         D => BU25_D,
         C => BU25_C,
         CE => BU25_CE,
         Q => BU25_Q
      );

   BU26_D <= n170;
   BU26_CE <= n180;
   BU26_CLK <= n183;
   BU26_A0 <= '0';
   BU26_A1 <= '1';
   BU26_A2 <= '0';
   BU26_A3 <= '0';
   n959 <= BU26_Q;
   BU26 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU26_D,
         CE => BU26_CE,
         CLK => BU26_CLK,
         A0 => BU26_A0,
         A1 => BU26_A1,
         A2 => BU26_A2,
         A3 => BU26_A3,
         Q => BU26_Q
      );

   BU28_D <= n959;
   BU28_C <= n183;
   BU28_CE <= n180;
   n614 <= BU28_Q;
   BU28 : FDE
      PORT MAP (
         D => BU28_D,
         C => BU28_C,
         CE => BU28_CE,
         Q => BU28_Q
      );

   BU29_D <= n171;
   BU29_CE <= n180;
   BU29_CLK <= n183;
   BU29_A0 <= '0';
   BU29_A1 <= '1';
   BU29_A2 <= '0';
   BU29_A3 <= '0';
   n960 <= BU29_Q;
   BU29 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU29_D,
         CE => BU29_CE,
         CLK => BU29_CLK,
         A0 => BU29_A0,
         A1 => BU29_A1,
         A2 => BU29_A2,
         A3 => BU29_A3,
         Q => BU29_Q
      );

   BU31_D <= n960;
   BU31_C <= n183;
   BU31_CE <= n180;
   n613 <= BU31_Q;
   BU31 : FDE
      PORT MAP (
         D => BU31_D,
         C => BU31_C,
         CE => BU31_CE,
         Q => BU31_Q
      );

   BU32_D <= n172;
   BU32_CE <= n180;
   BU32_CLK <= n183;
   BU32_A0 <= '0';
   BU32_A1 <= '1';
   BU32_A2 <= '0';
   BU32_A3 <= '0';
   n961 <= BU32_Q;
   BU32 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU32_D,
         CE => BU32_CE,
         CLK => BU32_CLK,
         A0 => BU32_A0,
         A1 => BU32_A1,
         A2 => BU32_A2,
         A3 => BU32_A3,
         Q => BU32_Q
      );

   BU34_D <= n961;
   BU34_C <= n183;
   BU34_CE <= n180;
   n612 <= BU34_Q;
   BU34 : FDE
      PORT MAP (
         D => BU34_D,
         C => BU34_C,
         CE => BU34_CE,
         Q => BU34_Q
      );

   BU35_D <= n173;
   BU35_CE <= n180;
   BU35_CLK <= n183;
   BU35_A0 <= '0';
   BU35_A1 <= '1';
   BU35_A2 <= '0';
   BU35_A3 <= '0';
   n962 <= BU35_Q;
   BU35 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU35_D,
         CE => BU35_CE,
         CLK => BU35_CLK,
         A0 => BU35_A0,
         A1 => BU35_A1,
         A2 => BU35_A2,
         A3 => BU35_A3,
         Q => BU35_Q
      );

   BU37_D <= n962;
   BU37_C <= n183;
   BU37_CE <= n180;
   n611 <= BU37_Q;
   BU37 : FDE
      PORT MAP (
         D => BU37_D,
         C => BU37_C,
         CE => BU37_CE,
         Q => BU37_Q
      );

   BU38_D <= n174;
   BU38_CE <= n180;
   BU38_CLK <= n183;
   BU38_A0 <= '0';
   BU38_A1 <= '1';
   BU38_A2 <= '0';
   BU38_A3 <= '0';
   n963 <= BU38_Q;
   BU38 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU38_D,
         CE => BU38_CE,
         CLK => BU38_CLK,
         A0 => BU38_A0,
         A1 => BU38_A1,
         A2 => BU38_A2,
         A3 => BU38_A3,
         Q => BU38_Q
      );

   BU40_D <= n963;
   BU40_C <= n183;
   BU40_CE <= n180;
   n610 <= BU40_Q;
   BU40 : FDE
      PORT MAP (
         D => BU40_D,
         C => BU40_C,
         CE => BU40_CE,
         Q => BU40_Q
      );

   BU41_D <= n175;
   BU41_CE <= n180;
   BU41_CLK <= n183;
   BU41_A0 <= '0';
   BU41_A1 <= '1';
   BU41_A2 <= '0';
   BU41_A3 <= '0';
   n964 <= BU41_Q;
   BU41 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU41_D,
         CE => BU41_CE,
         CLK => BU41_CLK,
         A0 => BU41_A0,
         A1 => BU41_A1,
         A2 => BU41_A2,
         A3 => BU41_A3,
         Q => BU41_Q
      );

   BU43_D <= n964;
   BU43_C <= n183;
   BU43_CE <= n180;
   n609 <= BU43_Q;
   BU43 : FDE
      PORT MAP (
         D => BU43_D,
         C => BU43_C,
         CE => BU43_CE,
         Q => BU43_Q
      );

   BU44_D <= n176;
   BU44_CE <= n180;
   BU44_CLK <= n183;
   BU44_A0 <= '0';
   BU44_A1 <= '1';
   BU44_A2 <= '0';
   BU44_A3 <= '0';
   n965 <= BU44_Q;
   BU44 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU44_D,
         CE => BU44_CE,
         CLK => BU44_CLK,
         A0 => BU44_A0,
         A1 => BU44_A1,
         A2 => BU44_A2,
         A3 => BU44_A3,
         Q => BU44_Q
      );

   BU46_D <= n965;
   BU46_C <= n183;
   BU46_CE <= n180;
   n608 <= BU46_Q;
   BU46 : FDE
      PORT MAP (
         D => BU46_D,
         C => BU46_C,
         CE => BU46_CE,
         Q => BU46_Q
      );

   BU47_D <= n177;
   BU47_CE <= n180;
   BU47_CLK <= n183;
   BU47_A0 <= '0';
   BU47_A1 <= '1';
   BU47_A2 <= '0';
   BU47_A3 <= '0';
   n966 <= BU47_Q;
   BU47 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU47_D,
         CE => BU47_CE,
         CLK => BU47_CLK,
         A0 => BU47_A0,
         A1 => BU47_A1,
         A2 => BU47_A2,
         A3 => BU47_A3,
         Q => BU47_Q
      );

   BU49_D <= n966;
   BU49_C <= n183;
   BU49_CE <= n180;
   n607 <= BU49_Q;
   BU49 : FDE
      PORT MAP (
         D => BU49_D,
         C => BU49_C,
         CE => BU49_CE,
         Q => BU49_Q
      );

   BU50_D <= n178;
   BU50_CE <= n180;
   BU50_CLK <= n183;
   BU50_A0 <= '0';
   BU50_A1 <= '1';
   BU50_A2 <= '0';
   BU50_A3 <= '0';
   n967 <= BU50_Q;
   BU50 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU50_D,
         CE => BU50_CE,
         CLK => BU50_CLK,
         A0 => BU50_A0,
         A1 => BU50_A1,
         A2 => BU50_A2,
         A3 => BU50_A3,
         Q => BU50_Q
      );

   BU52_D <= n967;
   BU52_C <= n183;
   BU52_CE <= n180;
   n606 <= BU52_Q;
   BU52 : FDE
      PORT MAP (
         D => BU52_D,
         C => BU52_C,
         CE => BU52_CE,
         Q => BU52_Q
      );

   BU53_D <= n179;
   BU53_CE <= n180;
   BU53_CLK <= n183;
   BU53_A0 <= '0';
   BU53_A1 <= '1';
   BU53_A2 <= '0';
   BU53_A3 <= '0';
   n968 <= BU53_Q;
   BU53 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU53_D,
         CE => BU53_CE,
         CLK => BU53_CLK,
         A0 => BU53_A0,
         A1 => BU53_A1,
         A2 => BU53_A2,
         A3 => BU53_A3,
         Q => BU53_Q
      );

   BU55_D <= n968;
   BU55_C <= n183;
   BU55_CE <= n180;
   n605 <= BU55_Q;
   BU55 : FDE
      PORT MAP (
         D => BU55_D,
         C => BU55_C,
         CE => BU55_CE,
         Q => BU55_Q
      );

   BU57_DATA(0) <= n189;
   BU57_DATA(1) <= n190;
   BU57_DATA(2) <= n191;
   BU57_DATA(3) <= n192;
   BU57_DATA(4) <= n193;
   BU57_DATA(5) <= n194;
   BU57_DATA(6) <= n195;
   BU57_DATA(7) <= n196;
   BU57_DATA(8) <= n197;
   BU57_DATA(9) <= n198;
   BU57_DATA(10) <= n199;
   BU57_DATA(11) <= n200;
   BU57_DATA(12) <= n201;
   BU57_DATA(13) <= n202;
   BU57_DATA(14) <= n203;
   BU57_DATA(15) <= n204;
   BU57_DATA(16) <= n205;
   BU57_DATA(17) <= n206;
   BU57_DATA(18) <= n207;
   BU57_DATA(19) <= n208;
   BU57_DATA(20) <= n209;
   BU57_DATA(21) <= n210;
   BU57_DATA(22) <= n211;
   BU57_DATA(23) <= n212;
   BU57_DATA(24) <= n213;
   BU57_DATA(25) <= n214;
   BU57_DATA(26) <= n215;
   BU57_DATA(27) <= n216;
   BU57_DATA(28) <= n217;
   BU57_DATA(29) <= n218;
   BU57_DATA(30) <= n219;
   BU57_DATA(31) <= n220;
   BU57_WE <= n322;
   BU57_CLK <= n183;
   BU57_CE <= n180;
   n370 <= BU57_RDY;
   n457 <= BU57_SINE(0);
   n456 <= BU57_SINE(1);
   n455 <= BU57_SINE(2);
   n454 <= BU57_SINE(3);
   n453 <= BU57_SINE(4);
   n452 <= BU57_SINE(5);
   n451 <= BU57_SINE(6);
   n450 <= BU57_SINE(7);
   n449 <= BU57_SINE(8);
   n448 <= BU57_SINE(9);
   n447 <= BU57_SINE(10);
   n446 <= BU57_SINE(11);
   n445 <= BU57_SINE(12);
   n444 <= BU57_SINE(13);
   n443 <= BU57_SINE(14);
   n661 <= BU57_COSINE(0);
   n660 <= BU57_COSINE(1);
   n659 <= BU57_COSINE(2);
   n658 <= BU57_COSINE(3);
   n657 <= BU57_COSINE(4);
   n656 <= BU57_COSINE(5);
   n655 <= BU57_COSINE(6);
   n654 <= BU57_COSINE(7);
   n653 <= BU57_COSINE(8);
   n652 <= BU57_COSINE(9);
   n651 <= BU57_COSINE(10);
   n650 <= BU57_COSINE(11);
   n649 <= BU57_COSINE(12);
   n648 <= BU57_COSINE(13);
   n647 <= BU57_COSINE(14);
   BU57 : C_DDS_V4_1
      GENERIC MAP (
         c_phase_offset_value => "00000000000000000000000000000000",
         c_phase_increment_value => "01001100110011001100110011001101",
         c_has_rdy => 1,
         c_has_sclr => 0,
         c_phase_offset => 0,
         c_data_width => 32,
         c_accumulator_latency => 1,
         c_enable_rlocs => 0,
         c_phase_angle_width => 13,
         c_has_rfd => 0,
         c_phase_increment => 1,
         c_negative_sine => 0,
         c_latency => 4,
         c_has_ce => 1,
         c_has_aclr => 0,
         c_outputs_required => 2,
         c_pipelined => 1,
         c_accumulator_width => 32,
         c_mem_type => 1,
         c_negative_cosine => 0,
         c_noise_shaping => 1,
         c_output_width => 15
      )
      PORT MAP (
         DATA => BU57_DATA,
         WE => BU57_WE,
         CLK => BU57_CLK,
         CE => BU57_CE,
         RDY => BU57_RDY,
         SINE => BU57_SINE,
         COSINE => BU57_COSINE
      );

   BU1294_I0 <= n370;
   BU1294_I1 <= n371;
   BU1294_I2 <= '0';
   BU1294_I3 <= '0';
   n369 <= BU1294_O;
   BU1294 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU1294_I0,
         I1 => BU1294_I1,
         I2 => BU1294_I2,
         I3 => BU1294_I3,
         O => BU1294_O
      );

   BU1296_clk <= n183;
   BU1296_a(13) <= n605;
   BU1296_a(12) <= n606;
   BU1296_a(11) <= n607;
   BU1296_a(10) <= n608;
   BU1296_a(9) <= n609;
   BU1296_a(8) <= n610;
   BU1296_a(7) <= n611;
   BU1296_a(6) <= n612;
   BU1296_a(5) <= n613;
   BU1296_a(4) <= n614;
   BU1296_a(3) <= n615;
   BU1296_a(2) <= n616;
   BU1296_a(1) <= n617;
   BU1296_a(0) <= n618;
   BU1296_b(14) <= n443;
   BU1296_b(13) <= n444;
   BU1296_b(12) <= n445;
   BU1296_b(11) <= n446;
   BU1296_b(10) <= n447;
   BU1296_b(9) <= n448;
   BU1296_b(8) <= n449;
   BU1296_b(7) <= n450;
   BU1296_b(6) <= n451;
   BU1296_b(5) <= n452;
   BU1296_b(4) <= n453;
   BU1296_b(3) <= n454;
   BU1296_b(2) <= n455;
   BU1296_b(1) <= n456;
   BU1296_b(0) <= n457;
   n488 <= BU1296_q(28);
   n489 <= BU1296_q(27);
   n490 <= BU1296_q(26);
   n491 <= BU1296_q(25);
   n492 <= BU1296_q(24);
   n493 <= BU1296_q(23);
   n494 <= BU1296_q(22);
   n495 <= BU1296_q(21);
   n496 <= BU1296_q(20);
   n497 <= BU1296_q(19);
   n498 <= BU1296_q(18);
   n499 <= BU1296_q(17);
   n500 <= BU1296_q(16);
   n501 <= BU1296_q(15);
   n502 <= BU1296_q(14);
   n503 <= BU1296_q(13);
   n504 <= BU1296_q(12);
   n505 <= BU1296_q(11);
   n506 <= BU1296_q(10);
   n507 <= BU1296_q(9);
   n508 <= BU1296_q(8);
   n509 <= BU1296_q(7);
   n510 <= BU1296_q(6);
   n511 <= BU1296_q(5);
   n512 <= BU1296_q(4);
   n513 <= BU1296_q(3);
   n514 <= BU1296_q(2);
   n515 <= BU1296_q(1);
   n516 <= BU1296_q(0);
   BU1296_a_signed <= '0';
   BU1296_loadb <= '0';
   BU1296_swapb <= '0';
   BU1296_ce <= '1';
   BU1296_aclr <= '0';
   BU1296_sclr <= '0';
   BU1296_nd <= n369;
   n575 <= BU1296_rdy;
   BU1296 : mult_gen_v5_0
      GENERIC MAP (
         c_a_width => 14,
         c_out_width => 29,
         c_b_type => 0,
         c_has_b => 1,
         c_has_rdy => 1,
         bram_addr_width => 8,
         c_has_sclr => 0,
         c_has_nd => 1,
         c_reg_a_b_inputs => 1,
         c_enable_rlocs => 0,
         c_has_rfd => 1,
         c_mult_type => 1,
         c_has_swapb => 0,
         c_baat => 14,
         c_use_luts => 1,
         c_has_load_done => 0,
         c_has_a_signed => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 1,
         c_output_hold => 0,
         c_stack_adders => 0,
         c_mem_type => 0,
         c_b_constant => 0,
         c_has_q => 1,
         c_has_loadb => 0,
         c_pipeline => 1,
         c_has_o => 0,
         c_standalone => 1,
         c_mem_init_prefix => "mem",
         c_a_type => 0,
         c_b_width => 15,
         c_sqm_type => 0,
         c_b_value => "0"
      )
      PORT MAP (
         clk => BU1296_clk,
         a => BU1296_a,
         b => BU1296_b,
         o => BU1296_o,
         q => BU1296_q,
         a_signed => BU1296_a_signed,
         loadb => BU1296_loadb,
         load_done => BU1296_load_done,
         swapb => BU1296_swapb,
         ce => BU1296_ce,
         aclr => BU1296_aclr,
         sclr => BU1296_sclr,
         rfd => BU1296_rfd,
         nd => BU1296_nd,
         rdy => BU1296_rdy
      );

   BU1517_I(0) <= n516;
   BU1517_I(1) <= n515;
   BU1517_I(2) <= n514;
   BU1517_I(3) <= n513;
   BU1517_I(4) <= n512;
   n1575 <= BU1517_O;
   BU1517 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 5,
         c_input_inv_mask => "01111"
      )
      PORT MAP (
         I => BU1517_I,
         O => BU1517_O
      );

   BU1526_I0 <= n511;
   BU1526_I1 <= n512;
   BU1526_I2 <= n1575;
   BU1526_I3 <= '0';
   n1572 <= BU1526_O;
   BU1526 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU1526_I0,
         I1 => BU1526_I1,
         I2 => BU1526_I2,
         I3 => BU1526_I3,
         O => BU1526_O
      );

   BU1527_A(0) <= n511;
   BU1527_A(1) <= n510;
   BU1527_A(2) <= n509;
   BU1527_A(3) <= n508;
   BU1527_A(4) <= n507;
   BU1527_A(5) <= n506;
   BU1527_A(6) <= n505;
   BU1527_A(7) <= n504;
   BU1527_A(8) <= n503;
   BU1527_A(9) <= n502;
   BU1527_A(10) <= n501;
   BU1527_A(11) <= n500;
   BU1527_A(12) <= n499;
   BU1527_A(13) <= n498;
   BU1527_A(14) <= n497;
   BU1527_A(15) <= n496;
   BU1527_A(16) <= n495;
   BU1527_A(17) <= n494;
   BU1527_A(18) <= n493;
   BU1527_A(19) <= n492;
   BU1527_A(20) <= n491;
   BU1527_A(21) <= n490;
   BU1527_A(22) <= n489;
   BU1527_A(23) <= n488;
   BU1527_B(0) <= n1572;
   n1547 <= BU1527_S(0);
   n1548 <= BU1527_S(1);
   n1549 <= BU1527_S(2);
   n1550 <= BU1527_S(3);
   n1551 <= BU1527_S(4);
   n1552 <= BU1527_S(5);
   n1553 <= BU1527_S(6);
   n1554 <= BU1527_S(7);
   n1555 <= BU1527_S(8);
   n1556 <= BU1527_S(9);
   n1557 <= BU1527_S(10);
   n1558 <= BU1527_S(11);
   n1559 <= BU1527_S(12);
   n1560 <= BU1527_S(13);
   n1561 <= BU1527_S(14);
   n1562 <= BU1527_S(15);
   n1563 <= BU1527_S(16);
   n1564 <= BU1527_S(17);
   n1565 <= BU1527_S(18);
   n1566 <= BU1527_S(19);
   n1567 <= BU1527_S(20);
   n1568 <= BU1527_S(21);
   n1569 <= BU1527_S(22);
   n1570 <= BU1527_S(23);
   BU1527 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU1527_A,
         B => BU1527_B,
         S => BU1527_S
      );

   BU1628_I0 <= n488;
   BU1628_I1 <= n489;
   BU1628_I2 <= n1570;
   BU1628_I3 <= '0';
   n1581 <= BU1628_O;
   BU1628 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU1628_I0,
         I1 => BU1628_I1,
         I2 => BU1628_I2,
         I3 => BU1628_I3,
         O => BU1628_O
      );

   BU1630_I0 <= n488;
   BU1630_I1 <= n1570;
   BU1630_I2 <= '0';
   BU1630_I3 <= '0';
   n1583 <= BU1630_O;
   BU1630 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU1630_I0,
         I1 => BU1630_I1,
         I2 => BU1630_I2,
         I3 => BU1630_I3,
         O => BU1630_O
      );

   BU1631_D(0) <= n1547;
   BU1631_D(1) <= n1548;
   BU1631_D(2) <= n1549;
   BU1631_D(3) <= n1550;
   BU1631_D(4) <= n1551;
   BU1631_D(5) <= n1552;
   BU1631_D(6) <= n1553;
   BU1631_D(7) <= n1554;
   BU1631_D(8) <= n1555;
   BU1631_D(9) <= n1556;
   BU1631_D(10) <= n1557;
   BU1631_D(11) <= n1558;
   BU1631_D(12) <= n1559;
   BU1631_D(13) <= n1560;
   BU1631_D(14) <= n1561;
   BU1631_D(15) <= n1562;
   BU1631_D(16) <= n1563;
   BU1631_D(17) <= n1564;
   BU1631_D(18) <= n1565;
   BU1631_D(19) <= n1566;
   BU1631_D(20) <= n1567;
   BU1631_D(21) <= n1568;
   BU1631_D(22) <= n1569;
   n3 <= BU1631_Q(0);
   n4 <= BU1631_Q(1);
   n5 <= BU1631_Q(2);
   n6 <= BU1631_Q(3);
   n7 <= BU1631_Q(4);
   n8 <= BU1631_Q(5);
   n9 <= BU1631_Q(6);
   n10 <= BU1631_Q(7);
   n11 <= BU1631_Q(8);
   n12 <= BU1631_Q(9);
   n13 <= BU1631_Q(10);
   n14 <= BU1631_Q(11);
   n15 <= BU1631_Q(12);
   n16 <= BU1631_Q(13);
   n17 <= BU1631_Q(14);
   n18 <= BU1631_Q(15);
   n19 <= BU1631_Q(16);
   n20 <= BU1631_Q(17);
   n21 <= BU1631_Q(18);
   n22 <= BU1631_Q(19);
   n23 <= BU1631_Q(20);
   n24 <= BU1631_Q(21);
   n25 <= BU1631_Q(22);
   BU1631_CLK <= n183;
   BU1631_SCLR <= n1581;
   BU1631_SSET <= n1583;
   BU1631 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU1631_D,
         Q => BU1631_Q,
         CLK => BU1631_CLK,
         SCLR => BU1631_SCLR,
         SSET => BU1631_SSET
      );

   BU1724_D(0) <= n1570;
   n26 <= BU1724_Q(0);
   BU1724_CLK <= n183;
   BU1724_SCLR <= n1583;
   BU1724_SSET <= n1581;
   BU1724 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU1724_D,
         Q => BU1724_Q,
         CLK => BU1724_CLK,
         SCLR => BU1724_SCLR,
         SSET => BU1724_SSET
      );

   BU1729_CLK <= n183;
   BU1729_D(0) <= n575;
   n2 <= BU1729_Q(0);
   BU1729 : C_SHIFT_RAM_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_read_mif => 0,
         c_has_a => 0,
         c_sync_priority => 0,
         c_has_sclr => 0,
         c_width => 1,
         c_enable_rlocs => 0,
         c_default_data_radix => 2,
         c_generate_mif => 0,
         c_ainit_val => "0",
         c_has_ce => 0,
         c_has_aclr => 0,
         c_mem_init_radix => 2,
         c_sync_enable => 0,
         c_depth => 1,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_shift_type => 0,
         c_mem_init_file => "null",
         c_default_data => "0",
         c_reg_last_bit => 1,
         c_addr_width => 0
      )
      PORT MAP (
         CLK => BU1729_CLK,
         D => BU1729_D,
         Q => BU1729_Q
      );

   BU1734_clk <= n183;
   BU1734_a(13) <= n605;
   BU1734_a(12) <= n606;
   BU1734_a(11) <= n607;
   BU1734_a(10) <= n608;
   BU1734_a(9) <= n609;
   BU1734_a(8) <= n610;
   BU1734_a(7) <= n611;
   BU1734_a(6) <= n612;
   BU1734_a(5) <= n613;
   BU1734_a(4) <= n614;
   BU1734_a(3) <= n615;
   BU1734_a(2) <= n616;
   BU1734_a(1) <= n617;
   BU1734_a(0) <= n618;
   BU1734_b(14) <= n647;
   BU1734_b(13) <= n648;
   BU1734_b(12) <= n649;
   BU1734_b(11) <= n650;
   BU1734_b(10) <= n651;
   BU1734_b(9) <= n652;
   BU1734_b(8) <= n653;
   BU1734_b(7) <= n654;
   BU1734_b(6) <= n655;
   BU1734_b(5) <= n656;
   BU1734_b(4) <= n657;
   BU1734_b(3) <= n658;
   BU1734_b(2) <= n659;
   BU1734_b(1) <= n660;
   BU1734_b(0) <= n661;
   n692 <= BU1734_q(28);
   n693 <= BU1734_q(27);
   n694 <= BU1734_q(26);
   n695 <= BU1734_q(25);
   n696 <= BU1734_q(24);
   n697 <= BU1734_q(23);
   n698 <= BU1734_q(22);
   n699 <= BU1734_q(21);
   n700 <= BU1734_q(20);
   n701 <= BU1734_q(19);
   n702 <= BU1734_q(18);
   n703 <= BU1734_q(17);
   n704 <= BU1734_q(16);
   n705 <= BU1734_q(15);
   n706 <= BU1734_q(14);
   n707 <= BU1734_q(13);
   n708 <= BU1734_q(12);
   n709 <= BU1734_q(11);
   n710 <= BU1734_q(10);
   n711 <= BU1734_q(9);
   n712 <= BU1734_q(8);
   n713 <= BU1734_q(7);
   n714 <= BU1734_q(6);
   n715 <= BU1734_q(5);
   n716 <= BU1734_q(4);
   n717 <= BU1734_q(3);
   n718 <= BU1734_q(2);
   n719 <= BU1734_q(1);
   n720 <= BU1734_q(0);
   BU1734_a_signed <= '0';
   BU1734_loadb <= '0';
   BU1734_swapb <= '0';
   BU1734_ce <= '1';
   BU1734_aclr <= '0';
   BU1734_sclr <= '0';
   BU1734_nd <= n369;
   BU1734 : mult_gen_v5_0
      GENERIC MAP (
         c_a_width => 14,
         c_out_width => 29,
         c_b_type => 0,
         c_has_b => 1,
         c_has_rdy => 1,
         bram_addr_width => 8,
         c_has_sclr => 0,
         c_has_nd => 1,
         c_reg_a_b_inputs => 1,
         c_enable_rlocs => 0,
         c_has_rfd => 1,
         c_mult_type => 1,
         c_has_swapb => 0,
         c_baat => 14,
         c_use_luts => 1,
         c_has_load_done => 0,
         c_has_a_signed => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 1,
         c_output_hold => 0,
         c_stack_adders => 0,
         c_mem_type => 0,
         c_b_constant => 0,
         c_has_q => 1,
         c_has_loadb => 0,
         c_pipeline => 1,
         c_has_o => 0,
         c_standalone => 1,
         c_mem_init_prefix => "mem",
         c_a_type => 0,
         c_b_width => 15,
         c_sqm_type => 0,
         c_b_value => "0"
      )
      PORT MAP (
         clk => BU1734_clk,
         a => BU1734_a,
         b => BU1734_b,
         o => BU1734_o,
         q => BU1734_q,
         a_signed => BU1734_a_signed,
         loadb => BU1734_loadb,
         load_done => BU1734_load_done,
         swapb => BU1734_swapb,
         ce => BU1734_ce,
         aclr => BU1734_aclr,
         sclr => BU1734_sclr,
         rfd => BU1734_rfd,
         nd => BU1734_nd,
         rdy => BU1734_rdy
      );

   BU1955_I(0) <= n720;
   BU1955_I(1) <= n719;
   BU1955_I(2) <= n718;
   BU1955_I(3) <= n717;
   BU1955_I(4) <= n716;
   n2218 <= BU1955_O;
   BU1955 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 5,
         c_input_inv_mask => "01111"
      )
      PORT MAP (
         I => BU1955_I,
         O => BU1955_O
      );

   BU1964_I0 <= n715;
   BU1964_I1 <= n716;
   BU1964_I2 <= n2218;
   BU1964_I3 <= '0';
   n2215 <= BU1964_O;
   BU1964 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU1964_I0,
         I1 => BU1964_I1,
         I2 => BU1964_I2,
         I3 => BU1964_I3,
         O => BU1964_O
      );

   BU1965_A(0) <= n715;
   BU1965_A(1) <= n714;
   BU1965_A(2) <= n713;
   BU1965_A(3) <= n712;
   BU1965_A(4) <= n711;
   BU1965_A(5) <= n710;
   BU1965_A(6) <= n709;
   BU1965_A(7) <= n708;
   BU1965_A(8) <= n707;
   BU1965_A(9) <= n706;
   BU1965_A(10) <= n705;
   BU1965_A(11) <= n704;
   BU1965_A(12) <= n703;
   BU1965_A(13) <= n702;
   BU1965_A(14) <= n701;
   BU1965_A(15) <= n700;
   BU1965_A(16) <= n699;
   BU1965_A(17) <= n698;
   BU1965_A(18) <= n697;
   BU1965_A(19) <= n696;
   BU1965_A(20) <= n695;
   BU1965_A(21) <= n694;
   BU1965_A(22) <= n693;
   BU1965_A(23) <= n692;
   BU1965_B(0) <= n2215;
   n2190 <= BU1965_S(0);
   n2191 <= BU1965_S(1);
   n2192 <= BU1965_S(2);
   n2193 <= BU1965_S(3);
   n2194 <= BU1965_S(4);
   n2195 <= BU1965_S(5);
   n2196 <= BU1965_S(6);
   n2197 <= BU1965_S(7);
   n2198 <= BU1965_S(8);
   n2199 <= BU1965_S(9);
   n2200 <= BU1965_S(10);
   n2201 <= BU1965_S(11);
   n2202 <= BU1965_S(12);
   n2203 <= BU1965_S(13);
   n2204 <= BU1965_S(14);
   n2205 <= BU1965_S(15);
   n2206 <= BU1965_S(16);
   n2207 <= BU1965_S(17);
   n2208 <= BU1965_S(18);
   n2209 <= BU1965_S(19);
   n2210 <= BU1965_S(20);
   n2211 <= BU1965_S(21);
   n2212 <= BU1965_S(22);
   n2213 <= BU1965_S(23);
   BU1965 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU1965_A,
         B => BU1965_B,
         S => BU1965_S
      );

   BU2066_I0 <= n692;
   BU2066_I1 <= n693;
   BU2066_I2 <= n2213;
   BU2066_I3 <= '0';
   n2224 <= BU2066_O;
   BU2066 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU2066_I0,
         I1 => BU2066_I1,
         I2 => BU2066_I2,
         I3 => BU2066_I3,
         O => BU2066_O
      );

   BU2068_I0 <= n692;
   BU2068_I1 <= n2213;
   BU2068_I2 <= '0';
   BU2068_I3 <= '0';
   n2226 <= BU2068_O;
   BU2068 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU2068_I0,
         I1 => BU2068_I1,
         I2 => BU2068_I2,
         I3 => BU2068_I3,
         O => BU2068_O
      );

   BU2069_D(0) <= n2190;
   BU2069_D(1) <= n2191;
   BU2069_D(2) <= n2192;
   BU2069_D(3) <= n2193;
   BU2069_D(4) <= n2194;
   BU2069_D(5) <= n2195;
   BU2069_D(6) <= n2196;
   BU2069_D(7) <= n2197;
   BU2069_D(8) <= n2198;
   BU2069_D(9) <= n2199;
   BU2069_D(10) <= n2200;
   BU2069_D(11) <= n2201;
   BU2069_D(12) <= n2202;
   BU2069_D(13) <= n2203;
   BU2069_D(14) <= n2204;
   BU2069_D(15) <= n2205;
   BU2069_D(16) <= n2206;
   BU2069_D(17) <= n2207;
   BU2069_D(18) <= n2208;
   BU2069_D(19) <= n2209;
   BU2069_D(20) <= n2210;
   BU2069_D(21) <= n2211;
   BU2069_D(22) <= n2212;
   n27 <= BU2069_Q(0);
   n28 <= BU2069_Q(1);
   n29 <= BU2069_Q(2);
   n30 <= BU2069_Q(3);
   n31 <= BU2069_Q(4);
   n32 <= BU2069_Q(5);
   n33 <= BU2069_Q(6);
   n34 <= BU2069_Q(7);
   n35 <= BU2069_Q(8);
   n36 <= BU2069_Q(9);
   n37 <= BU2069_Q(10);
   n38 <= BU2069_Q(11);
   n39 <= BU2069_Q(12);
   n40 <= BU2069_Q(13);
   n41 <= BU2069_Q(14);
   n42 <= BU2069_Q(15);
   n43 <= BU2069_Q(16);
   n44 <= BU2069_Q(17);
   n45 <= BU2069_Q(18);
   n46 <= BU2069_Q(19);
   n47 <= BU2069_Q(20);
   n48 <= BU2069_Q(21);
   n49 <= BU2069_Q(22);
   BU2069_CLK <= n183;
   BU2069_SCLR <= n2224;
   BU2069_SSET <= n2226;
   BU2069 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2069_D,
         Q => BU2069_Q,
         CLK => BU2069_CLK,
         SCLR => BU2069_SCLR,
         SSET => BU2069_SSET
      );

   BU2162_D(0) <= n2213;
   n50 <= BU2162_Q(0);
   BU2162_CLK <= n183;
   BU2162_SCLR <= n2226;
   BU2162_SSET <= n2224;
   BU2162 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2162_D,
         Q => BU2162_Q,
         CLK => BU2162_CLK,
         SCLR => BU2162_SCLR,
         SSET => BU2162_SSET
      );

   BU2457_D <= n2754;
   BU2457_C <= n183;
   BU2457_CE <= '1';
   n2705 <= BU2457_Q;
   BU2457 : FDE
      PORT MAP (
         D => BU2457_D,
         C => BU2457_C,
         CE => BU2457_CE,
         Q => BU2457_Q
      );

   BU2461_I(0) <= n2707;
   BU2461_I(1) <= n2708;
   BU2461_I(2) <= n2709;
   BU2461_I(3) <= n2710;
   BU2461_I(4) <= n2711;
   BU2461_I(5) <= n2712;
   BU2461_I(6) <= n2713;
   BU2461_I(7) <= n2714;
   BU2461_I(8) <= n2715;
   BU2461_I(9) <= n2716;
   BU2461_I(10) <= n2717;
   BU2461_I(11) <= n2718;
   BU2461_I(12) <= n2719;
   BU2461_I(13) <= n2720;
   BU2461_I(14) <= n2721;
   BU2461_I(15) <= n2722;
   BU2461_I(16) <= n2723;
   BU2461_I(17) <= n2724;
   BU2461_I(18) <= n2725;
   BU2461_I(19) <= n2726;
   BU2461_I(20) <= n2727;
   BU2461_I(21) <= n2728;
   BU2461_I(22) <= n2729;
   n3070 <= BU2461_O;
   BU2461 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 23,
         c_input_inv_mask => "01111111111111111111111"
      )
      PORT MAP (
         I => BU2461_I,
         O => BU2461_O
      );

   BU2489_I0 <= n2730;
   BU2489_I1 <= n2729;
   BU2489_I2 <= n3070;
   BU2489_I3 <= '0';
   n3067 <= BU2489_O;
   BU2489 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU2489_I0,
         I1 => BU2489_I1,
         I2 => BU2489_I2,
         I3 => BU2489_I3,
         O => BU2489_O
      );

   BU2490_A(0) <= n2730;
   BU2490_A(1) <= n2731;
   BU2490_A(2) <= n2732;
   BU2490_A(3) <= n2733;
   BU2490_A(4) <= n2734;
   BU2490_A(5) <= n2735;
   BU2490_A(6) <= n2736;
   BU2490_A(7) <= n2737;
   BU2490_A(8) <= n2738;
   BU2490_A(9) <= n2739;
   BU2490_A(10) <= n2740;
   BU2490_A(11) <= n2741;
   BU2490_A(12) <= n2742;
   BU2490_A(13) <= n2743;
   BU2490_A(14) <= n2744;
   BU2490_A(15) <= n2745;
   BU2490_A(16) <= n2746;
   BU2490_A(17) <= n2747;
   BU2490_A(18) <= n2748;
   BU2490_A(19) <= n2749;
   BU2490_A(20) <= n2750;
   BU2490_A(21) <= n2751;
   BU2490_A(22) <= n2752;
   BU2490_A(23) <= n2753;
   BU2490_B(0) <= n3067;
   n3042 <= BU2490_S(0);
   n3043 <= BU2490_S(1);
   n3044 <= BU2490_S(2);
   n3045 <= BU2490_S(3);
   n3046 <= BU2490_S(4);
   n3047 <= BU2490_S(5);
   n3048 <= BU2490_S(6);
   n3049 <= BU2490_S(7);
   n3050 <= BU2490_S(8);
   n3051 <= BU2490_S(9);
   n3052 <= BU2490_S(10);
   n3053 <= BU2490_S(11);
   n3054 <= BU2490_S(12);
   n3055 <= BU2490_S(13);
   n3056 <= BU2490_S(14);
   n3057 <= BU2490_S(15);
   n3058 <= BU2490_S(16);
   n3059 <= BU2490_S(17);
   n3060 <= BU2490_S(18);
   n3061 <= BU2490_S(19);
   n3062 <= BU2490_S(20);
   n3063 <= BU2490_S(21);
   n3064 <= BU2490_S(22);
   n3065 <= BU2490_S(23);
   BU2490 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU2490_A,
         B => BU2490_B,
         S => BU2490_S
      );

   BU2591_I0 <= n2753;
   BU2591_I1 <= n2752;
   BU2591_I2 <= n3065;
   BU2591_I3 <= '0';
   n3094 <= BU2591_O;
   BU2591 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU2591_I0,
         I1 => BU2591_I1,
         I2 => BU2591_I2,
         I3 => BU2591_I3,
         O => BU2591_O
      );

   BU2593_I0 <= n2753;
   BU2593_I1 <= n3065;
   BU2593_I2 <= '0';
   BU2593_I3 <= '0';
   n3096 <= BU2593_O;
   BU2593 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU2593_I0,
         I1 => BU2593_I1,
         I2 => BU2593_I2,
         I3 => BU2593_I3,
         O => BU2593_O
      );

   BU2594_D(0) <= n3042;
   BU2594_D(1) <= n3043;
   BU2594_D(2) <= n3044;
   BU2594_D(3) <= n3045;
   BU2594_D(4) <= n3046;
   BU2594_D(5) <= n3047;
   BU2594_D(6) <= n3048;
   BU2594_D(7) <= n3049;
   BU2594_D(8) <= n3050;
   BU2594_D(9) <= n3051;
   BU2594_D(10) <= n3052;
   BU2594_D(11) <= n3053;
   BU2594_D(12) <= n3054;
   BU2594_D(13) <= n3055;
   BU2594_D(14) <= n3056;
   BU2594_D(15) <= n3057;
   BU2594_D(16) <= n3058;
   BU2594_D(17) <= n3059;
   BU2594_D(18) <= n3060;
   BU2594_D(19) <= n3061;
   BU2594_D(20) <= n3062;
   BU2594_D(21) <= n3063;
   BU2594_D(22) <= n3064;
   n2633 <= BU2594_Q(0);
   n2634 <= BU2594_Q(1);
   n2635 <= BU2594_Q(2);
   n2636 <= BU2594_Q(3);
   n2637 <= BU2594_Q(4);
   n2638 <= BU2594_Q(5);
   n2639 <= BU2594_Q(6);
   n2640 <= BU2594_Q(7);
   n2641 <= BU2594_Q(8);
   n2642 <= BU2594_Q(9);
   n2643 <= BU2594_Q(10);
   n2644 <= BU2594_Q(11);
   n2645 <= BU2594_Q(12);
   n2646 <= BU2594_Q(13);
   n2647 <= BU2594_Q(14);
   n2648 <= BU2594_Q(15);
   n2649 <= BU2594_Q(16);
   n2650 <= BU2594_Q(17);
   n2651 <= BU2594_Q(18);
   n2652 <= BU2594_Q(19);
   n2653 <= BU2594_Q(20);
   n2654 <= BU2594_Q(21);
   n2655 <= BU2594_Q(22);
   BU2594_CLK <= n183;
   BU2594_SCLR <= n3094;
   BU2594_SSET <= n3096;
   BU2594 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2594_D,
         Q => BU2594_Q,
         CLK => BU2594_CLK,
         SCLR => BU2594_SCLR,
         SSET => BU2594_SSET
      );

   BU2687_D(0) <= n3065;
   n2656 <= BU2687_Q(0);
   BU2687_CLK <= n183;
   BU2687_SCLR <= n3096;
   BU2687_SSET <= n3094;
   BU2687 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2687_D,
         Q => BU2687_Q,
         CLK => BU2687_CLK,
         SCLR => BU2687_SCLR,
         SSET => BU2687_SSET
      );

   BU7487_I(0) <= n2755;
   BU7487_I(1) <= n2756;
   BU7487_I(2) <= n2757;
   BU7487_I(3) <= n2758;
   BU7487_I(4) <= n2759;
   BU7487_I(5) <= n2760;
   BU7487_I(6) <= n2761;
   BU7487_I(7) <= n2762;
   BU7487_I(8) <= n2763;
   BU7487_I(9) <= n2764;
   BU7487_I(10) <= n2765;
   BU7487_I(11) <= n2766;
   BU7487_I(12) <= n2767;
   BU7487_I(13) <= n2768;
   BU7487_I(14) <= n2769;
   BU7487_I(15) <= n2770;
   BU7487_I(16) <= n2771;
   BU7487_I(17) <= n2772;
   BU7487_I(18) <= n2773;
   BU7487_I(19) <= n2774;
   BU7487_I(20) <= n2775;
   BU7487_I(21) <= n2776;
   BU7487_I(22) <= n2777;
   n3587 <= BU7487_O;
   BU7487 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 23,
         c_input_inv_mask => "01111111111111111111111"
      )
      PORT MAP (
         I => BU7487_I,
         O => BU7487_O
      );

   BU7515_I0 <= n2778;
   BU7515_I1 <= n2777;
   BU7515_I2 <= n3587;
   BU7515_I3 <= '0';
   n3584 <= BU7515_O;
   BU7515 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU7515_I0,
         I1 => BU7515_I1,
         I2 => BU7515_I2,
         I3 => BU7515_I3,
         O => BU7515_O
      );

   BU7516_A(0) <= n2778;
   BU7516_A(1) <= n2779;
   BU7516_A(2) <= n2780;
   BU7516_A(3) <= n2781;
   BU7516_A(4) <= n2782;
   BU7516_A(5) <= n2783;
   BU7516_A(6) <= n2784;
   BU7516_A(7) <= n2785;
   BU7516_A(8) <= n2786;
   BU7516_A(9) <= n2787;
   BU7516_A(10) <= n2788;
   BU7516_A(11) <= n2789;
   BU7516_A(12) <= n2790;
   BU7516_A(13) <= n2791;
   BU7516_A(14) <= n2792;
   BU7516_A(15) <= n2793;
   BU7516_A(16) <= n2794;
   BU7516_A(17) <= n2795;
   BU7516_A(18) <= n2796;
   BU7516_A(19) <= n2797;
   BU7516_A(20) <= n2798;
   BU7516_A(21) <= n2799;
   BU7516_A(22) <= n2800;
   BU7516_A(23) <= n2801;
   BU7516_B(0) <= n3584;
   n3559 <= BU7516_S(0);
   n3560 <= BU7516_S(1);
   n3561 <= BU7516_S(2);
   n3562 <= BU7516_S(3);
   n3563 <= BU7516_S(4);
   n3564 <= BU7516_S(5);
   n3565 <= BU7516_S(6);
   n3566 <= BU7516_S(7);
   n3567 <= BU7516_S(8);
   n3568 <= BU7516_S(9);
   n3569 <= BU7516_S(10);
   n3570 <= BU7516_S(11);
   n3571 <= BU7516_S(12);
   n3572 <= BU7516_S(13);
   n3573 <= BU7516_S(14);
   n3574 <= BU7516_S(15);
   n3575 <= BU7516_S(16);
   n3576 <= BU7516_S(17);
   n3577 <= BU7516_S(18);
   n3578 <= BU7516_S(19);
   n3579 <= BU7516_S(20);
   n3580 <= BU7516_S(21);
   n3581 <= BU7516_S(22);
   n3582 <= BU7516_S(23);
   BU7516 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU7516_A,
         B => BU7516_B,
         S => BU7516_S
      );

   BU7617_I0 <= n2801;
   BU7617_I1 <= n2800;
   BU7617_I2 <= n3582;
   BU7617_I3 <= '0';
   n3611 <= BU7617_O;
   BU7617 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU7617_I0,
         I1 => BU7617_I1,
         I2 => BU7617_I2,
         I3 => BU7617_I3,
         O => BU7617_O
      );

   BU7619_I0 <= n2801;
   BU7619_I1 <= n3582;
   BU7619_I2 <= '0';
   BU7619_I3 <= '0';
   n3613 <= BU7619_O;
   BU7619 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU7619_I0,
         I1 => BU7619_I1,
         I2 => BU7619_I2,
         I3 => BU7619_I3,
         O => BU7619_O
      );

   BU7620_D(0) <= n3559;
   BU7620_D(1) <= n3560;
   BU7620_D(2) <= n3561;
   BU7620_D(3) <= n3562;
   BU7620_D(4) <= n3563;
   BU7620_D(5) <= n3564;
   BU7620_D(6) <= n3565;
   BU7620_D(7) <= n3566;
   BU7620_D(8) <= n3567;
   BU7620_D(9) <= n3568;
   BU7620_D(10) <= n3569;
   BU7620_D(11) <= n3570;
   BU7620_D(12) <= n3571;
   BU7620_D(13) <= n3572;
   BU7620_D(14) <= n3573;
   BU7620_D(15) <= n3574;
   BU7620_D(16) <= n3575;
   BU7620_D(17) <= n3576;
   BU7620_D(18) <= n3577;
   BU7620_D(19) <= n3578;
   BU7620_D(20) <= n3579;
   BU7620_D(21) <= n3580;
   BU7620_D(22) <= n3581;
   n2657 <= BU7620_Q(0);
   n2658 <= BU7620_Q(1);
   n2659 <= BU7620_Q(2);
   n2660 <= BU7620_Q(3);
   n2661 <= BU7620_Q(4);
   n2662 <= BU7620_Q(5);
   n2663 <= BU7620_Q(6);
   n2664 <= BU7620_Q(7);
   n2665 <= BU7620_Q(8);
   n2666 <= BU7620_Q(9);
   n2667 <= BU7620_Q(10);
   n2668 <= BU7620_Q(11);
   n2669 <= BU7620_Q(12);
   n2670 <= BU7620_Q(13);
   n2671 <= BU7620_Q(14);
   n2672 <= BU7620_Q(15);
   n2673 <= BU7620_Q(16);
   n2674 <= BU7620_Q(17);
   n2675 <= BU7620_Q(18);
   n2676 <= BU7620_Q(19);
   n2677 <= BU7620_Q(20);
   n2678 <= BU7620_Q(21);
   n2679 <= BU7620_Q(22);
   BU7620_CLK <= n183;
   BU7620_SCLR <= n3611;
   BU7620_SSET <= n3613;
   BU7620 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU7620_D,
         Q => BU7620_Q,
         CLK => BU7620_CLK,
         SCLR => BU7620_SCLR,
         SSET => BU7620_SSET
      );

   BU7713_D(0) <= n3582;
   n2680 <= BU7713_Q(0);
   BU7713_CLK <= n183;
   BU7713_SCLR <= n3613;
   BU7713_SSET <= n3611;
   BU7713 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU7713_D,
         Q => BU7713_Q,
         CLK => BU7713_CLK,
         SCLR => BU7713_SCLR,
         SSET => BU7713_SSET
      );

   BU2173_D <= n2657;
   BU2173_C <= n183;
   BU2173_CE <= '1';
   n2681 <= BU2173_Q;
   BU2173 : FDE
      PORT MAP (
         D => BU2173_D,
         C => BU2173_C,
         CE => BU2173_CE,
         Q => BU2173_Q
      );

   BU2175_D <= n2658;
   BU2175_C <= n183;
   BU2175_CE <= '1';
   n2682 <= BU2175_Q;
   BU2175 : FDE
      PORT MAP (
         D => BU2175_D,
         C => BU2175_C,
         CE => BU2175_CE,
         Q => BU2175_Q
      );

   BU2177_D <= n2659;
   BU2177_C <= n183;
   BU2177_CE <= '1';
   n2683 <= BU2177_Q;
   BU2177 : FDE
      PORT MAP (
         D => BU2177_D,
         C => BU2177_C,
         CE => BU2177_CE,
         Q => BU2177_Q
      );

   BU2179_D <= n2660;
   BU2179_C <= n183;
   BU2179_CE <= '1';
   n2684 <= BU2179_Q;
   BU2179 : FDE
      PORT MAP (
         D => BU2179_D,
         C => BU2179_C,
         CE => BU2179_CE,
         Q => BU2179_Q
      );

   BU2181_D <= n2661;
   BU2181_C <= n183;
   BU2181_CE <= '1';
   n2685 <= BU2181_Q;
   BU2181 : FDE
      PORT MAP (
         D => BU2181_D,
         C => BU2181_C,
         CE => BU2181_CE,
         Q => BU2181_Q
      );

   BU2183_D <= n2662;
   BU2183_C <= n183;
   BU2183_CE <= '1';
   n2686 <= BU2183_Q;
   BU2183 : FDE
      PORT MAP (
         D => BU2183_D,
         C => BU2183_C,
         CE => BU2183_CE,
         Q => BU2183_Q
      );

   BU2185_D <= n2663;
   BU2185_C <= n183;
   BU2185_CE <= '1';
   n2687 <= BU2185_Q;
   BU2185 : FDE
      PORT MAP (
         D => BU2185_D,
         C => BU2185_C,
         CE => BU2185_CE,
         Q => BU2185_Q
      );

   BU2187_D <= n2664;
   BU2187_C <= n183;
   BU2187_CE <= '1';
   n2688 <= BU2187_Q;
   BU2187 : FDE
      PORT MAP (
         D => BU2187_D,
         C => BU2187_C,
         CE => BU2187_CE,
         Q => BU2187_Q
      );

   BU2189_D <= n2665;
   BU2189_C <= n183;
   BU2189_CE <= '1';
   n2689 <= BU2189_Q;
   BU2189 : FDE
      PORT MAP (
         D => BU2189_D,
         C => BU2189_C,
         CE => BU2189_CE,
         Q => BU2189_Q
      );

   BU2191_D <= n2666;
   BU2191_C <= n183;
   BU2191_CE <= '1';
   n2690 <= BU2191_Q;
   BU2191 : FDE
      PORT MAP (
         D => BU2191_D,
         C => BU2191_C,
         CE => BU2191_CE,
         Q => BU2191_Q
      );

   BU2193_D <= n2667;
   BU2193_C <= n183;
   BU2193_CE <= '1';
   n2691 <= BU2193_Q;
   BU2193 : FDE
      PORT MAP (
         D => BU2193_D,
         C => BU2193_C,
         CE => BU2193_CE,
         Q => BU2193_Q
      );

   BU2195_D <= n2668;
   BU2195_C <= n183;
   BU2195_CE <= '1';
   n2692 <= BU2195_Q;
   BU2195 : FDE
      PORT MAP (
         D => BU2195_D,
         C => BU2195_C,
         CE => BU2195_CE,
         Q => BU2195_Q
      );

   BU2197_D <= n2669;
   BU2197_C <= n183;
   BU2197_CE <= '1';
   n2693 <= BU2197_Q;
   BU2197 : FDE
      PORT MAP (
         D => BU2197_D,
         C => BU2197_C,
         CE => BU2197_CE,
         Q => BU2197_Q
      );

   BU2199_D <= n2670;
   BU2199_C <= n183;
   BU2199_CE <= '1';
   n2694 <= BU2199_Q;
   BU2199 : FDE
      PORT MAP (
         D => BU2199_D,
         C => BU2199_C,
         CE => BU2199_CE,
         Q => BU2199_Q
      );

   BU2201_D <= n2671;
   BU2201_C <= n183;
   BU2201_CE <= '1';
   n2695 <= BU2201_Q;
   BU2201 : FDE
      PORT MAP (
         D => BU2201_D,
         C => BU2201_C,
         CE => BU2201_CE,
         Q => BU2201_Q
      );

   BU2203_D <= n2672;
   BU2203_C <= n183;
   BU2203_CE <= '1';
   n2696 <= BU2203_Q;
   BU2203 : FDE
      PORT MAP (
         D => BU2203_D,
         C => BU2203_C,
         CE => BU2203_CE,
         Q => BU2203_Q
      );

   BU2205_D <= n2673;
   BU2205_C <= n183;
   BU2205_CE <= '1';
   n2697 <= BU2205_Q;
   BU2205 : FDE
      PORT MAP (
         D => BU2205_D,
         C => BU2205_C,
         CE => BU2205_CE,
         Q => BU2205_Q
      );

   BU2207_D <= n2674;
   BU2207_C <= n183;
   BU2207_CE <= '1';
   n2698 <= BU2207_Q;
   BU2207 : FDE
      PORT MAP (
         D => BU2207_D,
         C => BU2207_C,
         CE => BU2207_CE,
         Q => BU2207_Q
      );

   BU2209_D <= n2675;
   BU2209_C <= n183;
   BU2209_CE <= '1';
   n2699 <= BU2209_Q;
   BU2209 : FDE
      PORT MAP (
         D => BU2209_D,
         C => BU2209_C,
         CE => BU2209_CE,
         Q => BU2209_Q
      );

   BU2211_D <= n2676;
   BU2211_C <= n183;
   BU2211_CE <= '1';
   n2700 <= BU2211_Q;
   BU2211 : FDE
      PORT MAP (
         D => BU2211_D,
         C => BU2211_C,
         CE => BU2211_CE,
         Q => BU2211_Q
      );

   BU2213_D <= n2677;
   BU2213_C <= n183;
   BU2213_CE <= '1';
   n2701 <= BU2213_Q;
   BU2213 : FDE
      PORT MAP (
         D => BU2213_D,
         C => BU2213_C,
         CE => BU2213_CE,
         Q => BU2213_Q
      );

   BU2215_D <= n2678;
   BU2215_C <= n183;
   BU2215_CE <= '1';
   n2702 <= BU2215_Q;
   BU2215 : FDE
      PORT MAP (
         D => BU2215_D,
         C => BU2215_C,
         CE => BU2215_CE,
         Q => BU2215_Q
      );

   BU2217_D <= n2679;
   BU2217_C <= n183;
   BU2217_CE <= '1';
   n2703 <= BU2217_Q;
   BU2217 : FDE
      PORT MAP (
         D => BU2217_D,
         C => BU2217_C,
         CE => BU2217_CE,
         Q => BU2217_Q
      );

   BU2219_D <= n2680;
   BU2219_C <= n183;
   BU2219_CE <= '1';
   n2704 <= BU2219_Q;
   BU2219 : FDE
      PORT MAP (
         D => BU2219_D,
         C => BU2219_C,
         CE => BU2219_CE,
         Q => BU2219_Q
      );

   BU2220_MA(0) <= n2681;
   BU2220_MA(1) <= n2682;
   BU2220_MA(2) <= n2683;
   BU2220_MA(3) <= n2684;
   BU2220_MA(4) <= n2685;
   BU2220_MA(5) <= n2686;
   BU2220_MA(6) <= n2687;
   BU2220_MA(7) <= n2688;
   BU2220_MA(8) <= n2689;
   BU2220_MA(9) <= n2690;
   BU2220_MA(10) <= n2691;
   BU2220_MA(11) <= n2692;
   BU2220_MA(12) <= n2693;
   BU2220_MA(13) <= n2694;
   BU2220_MA(14) <= n2695;
   BU2220_MA(15) <= n2696;
   BU2220_MA(16) <= n2697;
   BU2220_MA(17) <= n2698;
   BU2220_MA(18) <= n2699;
   BU2220_MA(19) <= n2700;
   BU2220_MA(20) <= n2701;
   BU2220_MA(21) <= n2702;
   BU2220_MA(22) <= n2703;
   BU2220_MA(23) <= n2704;
   BU2220_MB(0) <= n2633;
   BU2220_MB(1) <= n2634;
   BU2220_MB(2) <= n2635;
   BU2220_MB(3) <= n2636;
   BU2220_MB(4) <= n2637;
   BU2220_MB(5) <= n2638;
   BU2220_MB(6) <= n2639;
   BU2220_MB(7) <= n2640;
   BU2220_MB(8) <= n2641;
   BU2220_MB(9) <= n2642;
   BU2220_MB(10) <= n2643;
   BU2220_MB(11) <= n2644;
   BU2220_MB(12) <= n2645;
   BU2220_MB(13) <= n2646;
   BU2220_MB(14) <= n2647;
   BU2220_MB(15) <= n2648;
   BU2220_MB(16) <= n2649;
   BU2220_MB(17) <= n2650;
   BU2220_MB(18) <= n2651;
   BU2220_MB(19) <= n2652;
   BU2220_MB(20) <= n2653;
   BU2220_MB(21) <= n2654;
   BU2220_MB(22) <= n2655;
   BU2220_MB(23) <= n2656;
   BU2220_S(0) <= n2705;
   n58 <= BU2220_Q(0);
   n59 <= BU2220_Q(1);
   n60 <= BU2220_Q(2);
   n61 <= BU2220_Q(3);
   n62 <= BU2220_Q(4);
   n63 <= BU2220_Q(5);
   n64 <= BU2220_Q(6);
   n65 <= BU2220_Q(7);
   n66 <= BU2220_Q(8);
   n67 <= BU2220_Q(9);
   n68 <= BU2220_Q(10);
   n69 <= BU2220_Q(11);
   n70 <= BU2220_Q(12);
   n71 <= BU2220_Q(13);
   n72 <= BU2220_Q(14);
   n73 <= BU2220_Q(15);
   n74 <= BU2220_Q(16);
   n75 <= BU2220_Q(17);
   n76 <= BU2220_Q(18);
   n77 <= BU2220_Q(19);
   n78 <= BU2220_Q(20);
   n79 <= BU2220_Q(21);
   n80 <= BU2220_Q(22);
   n81 <= BU2220_Q(23);
   BU2220_CLK <= n183;
   BU2220 : C_MUX_BUS_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_has_en => 0,
         c_sync_priority => 0,
         c_has_sclr => 0,
         c_width => 24,
         c_enable_rlocs => 0,
         c_sel_width => 1,
         c_latency => 1,
         c_ainit_val => "000000000000000000000000",
         c_has_ce => 0,
         c_mux_type => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "000000000000000000000000",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 1,
         c_has_o => 0,
         c_inputs => 2
      )
      PORT MAP (
         MA => BU2220_MA,
         MB => BU2220_MB,
         S => BU2220_S,
         Q => BU2220_Q,
         CLK => BU2220_CLK
      );

   BU2448_D <= n2705;
   BU2448_C <= n183;
   BU2448_CE <= '1';
   n2706 <= BU2448_Q;
   BU2448 : FDE
      PORT MAP (
         D => BU2448_D,
         C => BU2448_C,
         CE => BU2448_CE,
         Q => BU2448_Q
      );

   BU2452_I0 <= n2705;
   BU2452_I1 <= n2706;
   BU2452_I2 <= '0';
   BU2452_I3 <= '0';
   n4473 <= BU2452_O;
   BU2452 : LUT4
      GENERIC MAP (
         INIT  => X"eeee"
      )
      PORT MAP (
         I0 => BU2452_I0,
         I1 => BU2452_I1,
         I2 => BU2452_I2,
         I3 => BU2452_I3,
         O => BU2452_O
      );

   BU2453_D <= n4473;
   BU2453_C <= n183;
   BU2453_CE <= '1';
   n55 <= BU2453_Q;
   BU2453 : FDE
      PORT MAP (
         D => BU2453_D,
         C => BU2453_C,
         CE => BU2453_CE,
         Q => BU2453_Q
      );

   BU2692_DIN(0) <= n3;
   BU2692_DIN(1) <= n4;
   BU2692_DIN(2) <= n5;
   BU2692_DIN(3) <= n6;
   BU2692_DIN(4) <= n7;
   BU2692_DIN(5) <= n8;
   BU2692_DIN(6) <= n9;
   BU2692_DIN(7) <= n10;
   BU2692_DIN(8) <= n11;
   BU2692_DIN(9) <= n12;
   BU2692_DIN(10) <= n13;
   BU2692_DIN(11) <= n14;
   BU2692_DIN(12) <= n15;
   BU2692_DIN(13) <= n16;
   BU2692_DIN(14) <= n17;
   BU2692_DIN(15) <= n18;
   BU2692_DIN(16) <= n19;
   BU2692_DIN(17) <= n20;
   BU2692_DIN(18) <= n21;
   BU2692_DIN(19) <= n22;
   BU2692_DIN(20) <= n23;
   BU2692_DIN(21) <= n24;
   BU2692_DIN(22) <= n25;
   BU2692_DIN(23) <= n26;
   BU2692_ND <= n2;
   BU2692_CLK <= n183;
   n2707 <= BU2692_DOUT(0);
   n2708 <= BU2692_DOUT(1);
   n2709 <= BU2692_DOUT(2);
   n2710 <= BU2692_DOUT(3);
   n2711 <= BU2692_DOUT(4);
   n2712 <= BU2692_DOUT(5);
   n2713 <= BU2692_DOUT(6);
   n2714 <= BU2692_DOUT(7);
   n2715 <= BU2692_DOUT(8);
   n2716 <= BU2692_DOUT(9);
   n2717 <= BU2692_DOUT(10);
   n2718 <= BU2692_DOUT(11);
   n2719 <= BU2692_DOUT(12);
   n2720 <= BU2692_DOUT(13);
   n2721 <= BU2692_DOUT(14);
   n2722 <= BU2692_DOUT(15);
   n2723 <= BU2692_DOUT(16);
   n2724 <= BU2692_DOUT(17);
   n2725 <= BU2692_DOUT(18);
   n2726 <= BU2692_DOUT(19);
   n2727 <= BU2692_DOUT(20);
   n2728 <= BU2692_DOUT(21);
   n2729 <= BU2692_DOUT(22);
   n2730 <= BU2692_DOUT(23);
   n2731 <= BU2692_DOUT(24);
   n2732 <= BU2692_DOUT(25);
   n2733 <= BU2692_DOUT(26);
   n2734 <= BU2692_DOUT(27);
   n2735 <= BU2692_DOUT(28);
   n2736 <= BU2692_DOUT(29);
   n2737 <= BU2692_DOUT(30);
   n2738 <= BU2692_DOUT(31);
   n2739 <= BU2692_DOUT(32);
   n2740 <= BU2692_DOUT(33);
   n2741 <= BU2692_DOUT(34);
   n2742 <= BU2692_DOUT(35);
   n2743 <= BU2692_DOUT(36);
   n2744 <= BU2692_DOUT(37);
   n2745 <= BU2692_DOUT(38);
   n2746 <= BU2692_DOUT(39);
   n2747 <= BU2692_DOUT(40);
   n2748 <= BU2692_DOUT(41);
   n2749 <= BU2692_DOUT(42);
   n2750 <= BU2692_DOUT(43);
   n2751 <= BU2692_DOUT(44);
   n2752 <= BU2692_DOUT(45);
   n2753 <= BU2692_DOUT(46);
   n2754 <= BU2692_RDY;
   BU2692 : C_CIC_V3_0
      GENERIC MAP (
         c_differential_delay => 1,
         c_sample_rate_change_max => 16383,
         c_number_channels => 1,
         c_filter_type => 2,
         c_result_width => 47,
         c_enable_rlocs => 0,
         c_sample_rate_change => 10,
         c_latency => 1,
         c_sample_rate_change_min => 4,
         c_sample_rate_change_type => 2,
         c_data_width => 24,
         c_stages => 7
      )
      PORT MAP (
         DIN => BU2692_DIN,
         ND => BU2692_ND,
         RFD => BU2692_RFD,
         CLK => BU2692_CLK,
         DOUT => BU2692_DOUT,
         RDY => BU2692_RDY
      );

   BU7718_DIN(0) <= n27;
   BU7718_DIN(1) <= n28;
   BU7718_DIN(2) <= n29;
   BU7718_DIN(3) <= n30;
   BU7718_DIN(4) <= n31;
   BU7718_DIN(5) <= n32;
   BU7718_DIN(6) <= n33;
   BU7718_DIN(7) <= n34;
   BU7718_DIN(8) <= n35;
   BU7718_DIN(9) <= n36;
   BU7718_DIN(10) <= n37;
   BU7718_DIN(11) <= n38;
   BU7718_DIN(12) <= n39;
   BU7718_DIN(13) <= n40;
   BU7718_DIN(14) <= n41;
   BU7718_DIN(15) <= n42;
   BU7718_DIN(16) <= n43;
   BU7718_DIN(17) <= n44;
   BU7718_DIN(18) <= n45;
   BU7718_DIN(19) <= n46;
   BU7718_DIN(20) <= n47;
   BU7718_DIN(21) <= n48;
   BU7718_DIN(22) <= n49;
   BU7718_DIN(23) <= n50;
   BU7718_ND <= n2;
   BU7718_CLK <= n183;
   n2755 <= BU7718_DOUT(0);
   n2756 <= BU7718_DOUT(1);
   n2757 <= BU7718_DOUT(2);
   n2758 <= BU7718_DOUT(3);
   n2759 <= BU7718_DOUT(4);
   n2760 <= BU7718_DOUT(5);
   n2761 <= BU7718_DOUT(6);
   n2762 <= BU7718_DOUT(7);
   n2763 <= BU7718_DOUT(8);
   n2764 <= BU7718_DOUT(9);
   n2765 <= BU7718_DOUT(10);
   n2766 <= BU7718_DOUT(11);
   n2767 <= BU7718_DOUT(12);
   n2768 <= BU7718_DOUT(13);
   n2769 <= BU7718_DOUT(14);
   n2770 <= BU7718_DOUT(15);
   n2771 <= BU7718_DOUT(16);
   n2772 <= BU7718_DOUT(17);
   n2773 <= BU7718_DOUT(18);
   n2774 <= BU7718_DOUT(19);
   n2775 <= BU7718_DOUT(20);
   n2776 <= BU7718_DOUT(21);
   n2777 <= BU7718_DOUT(22);
   n2778 <= BU7718_DOUT(23);
   n2779 <= BU7718_DOUT(24);
   n2780 <= BU7718_DOUT(25);
   n2781 <= BU7718_DOUT(26);
   n2782 <= BU7718_DOUT(27);
   n2783 <= BU7718_DOUT(28);
   n2784 <= BU7718_DOUT(29);
   n2785 <= BU7718_DOUT(30);
   n2786 <= BU7718_DOUT(31);
   n2787 <= BU7718_DOUT(32);
   n2788 <= BU7718_DOUT(33);
   n2789 <= BU7718_DOUT(34);
   n2790 <= BU7718_DOUT(35);
   n2791 <= BU7718_DOUT(36);
   n2792 <= BU7718_DOUT(37);
   n2793 <= BU7718_DOUT(38);
   n2794 <= BU7718_DOUT(39);
   n2795 <= BU7718_DOUT(40);
   n2796 <= BU7718_DOUT(41);
   n2797 <= BU7718_DOUT(42);
   n2798 <= BU7718_DOUT(43);
   n2799 <= BU7718_DOUT(44);
   n2800 <= BU7718_DOUT(45);
   n2801 <= BU7718_DOUT(46);
   BU7718 : C_CIC_V3_0
      GENERIC MAP (
         c_differential_delay => 1,
         c_sample_rate_change_max => 16383,
         c_number_channels => 1,
         c_filter_type => 2,
         c_result_width => 47,
         c_enable_rlocs => 0,
         c_sample_rate_change => 10,
         c_latency => 1,
         c_sample_rate_change_min => 4,
         c_sample_rate_change_type => 2,
         c_data_width => 24,
         c_stages => 7
      )
      PORT MAP (
         DIN => BU7718_DIN,
         ND => BU7718_ND,
         RFD => BU7718_RFD,
         CLK => BU7718_CLK,
         DOUT => BU7718_DOUT,
         RDY => BU7718_RDY
      );

   BU12513_I0 <= n6747;
   BU12513_I1 <= n6719;
   BU12513_I2 <= '0';
   BU12513_I3 <= '0';
   n6746 <= BU12513_O;
   BU12513 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU12513_I0,
         I1 => BU12513_I1,
         I2 => BU12513_I2,
         I3 => BU12513_I3,
         O => BU12513_O
      );

   BU12518_I0 <= n55;
   BU12518_I1 <= '1';
   BU12518_I2 <= '0';
   BU12518_I3 <= '0';
   n6861 <= BU12518_O;
   BU12518 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU12518_I0,
         I1 => BU12518_I1,
         I2 => BU12518_I2,
         I3 => BU12518_I3,
         O => BU12518_O
      );

   BU12524_D <= '0';
   BU12524_CE <= n6861;
   BU12524_CLK <= n183;
   BU12524_A0 <= n6857;
   BU12524_A1 <= n6858;
   BU12524_A2 <= n6859;
   BU12524_A3 <= n6860;
   n6720 <= BU12524_Q;
   BU12524 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12524_D,
         CE => BU12524_CE,
         CLK => BU12524_CLK,
         A0 => BU12524_A0,
         A1 => BU12524_A1,
         A2 => BU12524_A2,
         A3 => BU12524_A3,
         Q => BU12524_Q
      );

   BU12525_D <= '0';
   BU12525_CE <= n6861;
   BU12525_CLK <= n183;
   BU12525_A0 <= n6857;
   BU12525_A1 <= n6858;
   BU12525_A2 <= n6859;
   BU12525_A3 <= n6860;
   n6721 <= BU12525_Q;
   BU12525 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12525_D,
         CE => BU12525_CE,
         CLK => BU12525_CLK,
         A0 => BU12525_A0,
         A1 => BU12525_A1,
         A2 => BU12525_A2,
         A3 => BU12525_A3,
         Q => BU12525_Q
      );

   BU12526_D <= n58;
   BU12526_CE <= n6861;
   BU12526_CLK <= n183;
   BU12526_A0 <= n6857;
   BU12526_A1 <= n6858;
   BU12526_A2 <= n6859;
   BU12526_A3 <= n6860;
   n6722 <= BU12526_Q;
   BU12526 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12526_D,
         CE => BU12526_CE,
         CLK => BU12526_CLK,
         A0 => BU12526_A0,
         A1 => BU12526_A1,
         A2 => BU12526_A2,
         A3 => BU12526_A3,
         Q => BU12526_Q
      );

   BU12527_D <= n59;
   BU12527_CE <= n6861;
   BU12527_CLK <= n183;
   BU12527_A0 <= n6857;
   BU12527_A1 <= n6858;
   BU12527_A2 <= n6859;
   BU12527_A3 <= n6860;
   n6723 <= BU12527_Q;
   BU12527 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12527_D,
         CE => BU12527_CE,
         CLK => BU12527_CLK,
         A0 => BU12527_A0,
         A1 => BU12527_A1,
         A2 => BU12527_A2,
         A3 => BU12527_A3,
         Q => BU12527_Q
      );

   BU12528_D <= n60;
   BU12528_CE <= n6861;
   BU12528_CLK <= n183;
   BU12528_A0 <= n6857;
   BU12528_A1 <= n6858;
   BU12528_A2 <= n6859;
   BU12528_A3 <= n6860;
   n6724 <= BU12528_Q;
   BU12528 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12528_D,
         CE => BU12528_CE,
         CLK => BU12528_CLK,
         A0 => BU12528_A0,
         A1 => BU12528_A1,
         A2 => BU12528_A2,
         A3 => BU12528_A3,
         Q => BU12528_Q
      );

   BU12529_D <= n61;
   BU12529_CE <= n6861;
   BU12529_CLK <= n183;
   BU12529_A0 <= n6857;
   BU12529_A1 <= n6858;
   BU12529_A2 <= n6859;
   BU12529_A3 <= n6860;
   n6725 <= BU12529_Q;
   BU12529 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12529_D,
         CE => BU12529_CE,
         CLK => BU12529_CLK,
         A0 => BU12529_A0,
         A1 => BU12529_A1,
         A2 => BU12529_A2,
         A3 => BU12529_A3,
         Q => BU12529_Q
      );

   BU12530_D <= n62;
   BU12530_CE <= n6861;
   BU12530_CLK <= n183;
   BU12530_A0 <= n6857;
   BU12530_A1 <= n6858;
   BU12530_A2 <= n6859;
   BU12530_A3 <= n6860;
   n6726 <= BU12530_Q;
   BU12530 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12530_D,
         CE => BU12530_CE,
         CLK => BU12530_CLK,
         A0 => BU12530_A0,
         A1 => BU12530_A1,
         A2 => BU12530_A2,
         A3 => BU12530_A3,
         Q => BU12530_Q
      );

   BU12531_D <= n63;
   BU12531_CE <= n6861;
   BU12531_CLK <= n183;
   BU12531_A0 <= n6857;
   BU12531_A1 <= n6858;
   BU12531_A2 <= n6859;
   BU12531_A3 <= n6860;
   n6727 <= BU12531_Q;
   BU12531 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12531_D,
         CE => BU12531_CE,
         CLK => BU12531_CLK,
         A0 => BU12531_A0,
         A1 => BU12531_A1,
         A2 => BU12531_A2,
         A3 => BU12531_A3,
         Q => BU12531_Q
      );

   BU12532_D <= n64;
   BU12532_CE <= n6861;
   BU12532_CLK <= n183;
   BU12532_A0 <= n6857;
   BU12532_A1 <= n6858;
   BU12532_A2 <= n6859;
   BU12532_A3 <= n6860;
   n6728 <= BU12532_Q;
   BU12532 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12532_D,
         CE => BU12532_CE,
         CLK => BU12532_CLK,
         A0 => BU12532_A0,
         A1 => BU12532_A1,
         A2 => BU12532_A2,
         A3 => BU12532_A3,
         Q => BU12532_Q
      );

   BU12533_D <= n65;
   BU12533_CE <= n6861;
   BU12533_CLK <= n183;
   BU12533_A0 <= n6857;
   BU12533_A1 <= n6858;
   BU12533_A2 <= n6859;
   BU12533_A3 <= n6860;
   n6729 <= BU12533_Q;
   BU12533 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12533_D,
         CE => BU12533_CE,
         CLK => BU12533_CLK,
         A0 => BU12533_A0,
         A1 => BU12533_A1,
         A2 => BU12533_A2,
         A3 => BU12533_A3,
         Q => BU12533_Q
      );

   BU12534_D <= n66;
   BU12534_CE <= n6861;
   BU12534_CLK <= n183;
   BU12534_A0 <= n6857;
   BU12534_A1 <= n6858;
   BU12534_A2 <= n6859;
   BU12534_A3 <= n6860;
   n6730 <= BU12534_Q;
   BU12534 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12534_D,
         CE => BU12534_CE,
         CLK => BU12534_CLK,
         A0 => BU12534_A0,
         A1 => BU12534_A1,
         A2 => BU12534_A2,
         A3 => BU12534_A3,
         Q => BU12534_Q
      );

   BU12535_D <= n67;
   BU12535_CE <= n6861;
   BU12535_CLK <= n183;
   BU12535_A0 <= n6857;
   BU12535_A1 <= n6858;
   BU12535_A2 <= n6859;
   BU12535_A3 <= n6860;
   n6731 <= BU12535_Q;
   BU12535 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12535_D,
         CE => BU12535_CE,
         CLK => BU12535_CLK,
         A0 => BU12535_A0,
         A1 => BU12535_A1,
         A2 => BU12535_A2,
         A3 => BU12535_A3,
         Q => BU12535_Q
      );

   BU12536_D <= n68;
   BU12536_CE <= n6861;
   BU12536_CLK <= n183;
   BU12536_A0 <= n6857;
   BU12536_A1 <= n6858;
   BU12536_A2 <= n6859;
   BU12536_A3 <= n6860;
   n6732 <= BU12536_Q;
   BU12536 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12536_D,
         CE => BU12536_CE,
         CLK => BU12536_CLK,
         A0 => BU12536_A0,
         A1 => BU12536_A1,
         A2 => BU12536_A2,
         A3 => BU12536_A3,
         Q => BU12536_Q
      );

   BU12537_D <= n69;
   BU12537_CE <= n6861;
   BU12537_CLK <= n183;
   BU12537_A0 <= n6857;
   BU12537_A1 <= n6858;
   BU12537_A2 <= n6859;
   BU12537_A3 <= n6860;
   n6733 <= BU12537_Q;
   BU12537 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12537_D,
         CE => BU12537_CE,
         CLK => BU12537_CLK,
         A0 => BU12537_A0,
         A1 => BU12537_A1,
         A2 => BU12537_A2,
         A3 => BU12537_A3,
         Q => BU12537_Q
      );

   BU12538_D <= n70;
   BU12538_CE <= n6861;
   BU12538_CLK <= n183;
   BU12538_A0 <= n6857;
   BU12538_A1 <= n6858;
   BU12538_A2 <= n6859;
   BU12538_A3 <= n6860;
   n6734 <= BU12538_Q;
   BU12538 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12538_D,
         CE => BU12538_CE,
         CLK => BU12538_CLK,
         A0 => BU12538_A0,
         A1 => BU12538_A1,
         A2 => BU12538_A2,
         A3 => BU12538_A3,
         Q => BU12538_Q
      );

   BU12539_D <= n71;
   BU12539_CE <= n6861;
   BU12539_CLK <= n183;
   BU12539_A0 <= n6857;
   BU12539_A1 <= n6858;
   BU12539_A2 <= n6859;
   BU12539_A3 <= n6860;
   n6735 <= BU12539_Q;
   BU12539 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12539_D,
         CE => BU12539_CE,
         CLK => BU12539_CLK,
         A0 => BU12539_A0,
         A1 => BU12539_A1,
         A2 => BU12539_A2,
         A3 => BU12539_A3,
         Q => BU12539_Q
      );

   BU12540_D <= n72;
   BU12540_CE <= n6861;
   BU12540_CLK <= n183;
   BU12540_A0 <= n6857;
   BU12540_A1 <= n6858;
   BU12540_A2 <= n6859;
   BU12540_A3 <= n6860;
   n6736 <= BU12540_Q;
   BU12540 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12540_D,
         CE => BU12540_CE,
         CLK => BU12540_CLK,
         A0 => BU12540_A0,
         A1 => BU12540_A1,
         A2 => BU12540_A2,
         A3 => BU12540_A3,
         Q => BU12540_Q
      );

   BU12541_D <= n73;
   BU12541_CE <= n6861;
   BU12541_CLK <= n183;
   BU12541_A0 <= n6857;
   BU12541_A1 <= n6858;
   BU12541_A2 <= n6859;
   BU12541_A3 <= n6860;
   n6737 <= BU12541_Q;
   BU12541 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12541_D,
         CE => BU12541_CE,
         CLK => BU12541_CLK,
         A0 => BU12541_A0,
         A1 => BU12541_A1,
         A2 => BU12541_A2,
         A3 => BU12541_A3,
         Q => BU12541_Q
      );

   BU12542_D <= n74;
   BU12542_CE <= n6861;
   BU12542_CLK <= n183;
   BU12542_A0 <= n6857;
   BU12542_A1 <= n6858;
   BU12542_A2 <= n6859;
   BU12542_A3 <= n6860;
   n6738 <= BU12542_Q;
   BU12542 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12542_D,
         CE => BU12542_CE,
         CLK => BU12542_CLK,
         A0 => BU12542_A0,
         A1 => BU12542_A1,
         A2 => BU12542_A2,
         A3 => BU12542_A3,
         Q => BU12542_Q
      );

   BU12543_D <= n75;
   BU12543_CE <= n6861;
   BU12543_CLK <= n183;
   BU12543_A0 <= n6857;
   BU12543_A1 <= n6858;
   BU12543_A2 <= n6859;
   BU12543_A3 <= n6860;
   n6739 <= BU12543_Q;
   BU12543 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12543_D,
         CE => BU12543_CE,
         CLK => BU12543_CLK,
         A0 => BU12543_A0,
         A1 => BU12543_A1,
         A2 => BU12543_A2,
         A3 => BU12543_A3,
         Q => BU12543_Q
      );

   BU12544_D <= n76;
   BU12544_CE <= n6861;
   BU12544_CLK <= n183;
   BU12544_A0 <= n6857;
   BU12544_A1 <= n6858;
   BU12544_A2 <= n6859;
   BU12544_A3 <= n6860;
   n6740 <= BU12544_Q;
   BU12544 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12544_D,
         CE => BU12544_CE,
         CLK => BU12544_CLK,
         A0 => BU12544_A0,
         A1 => BU12544_A1,
         A2 => BU12544_A2,
         A3 => BU12544_A3,
         Q => BU12544_Q
      );

   BU12545_D <= n77;
   BU12545_CE <= n6861;
   BU12545_CLK <= n183;
   BU12545_A0 <= n6857;
   BU12545_A1 <= n6858;
   BU12545_A2 <= n6859;
   BU12545_A3 <= n6860;
   n6741 <= BU12545_Q;
   BU12545 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12545_D,
         CE => BU12545_CE,
         CLK => BU12545_CLK,
         A0 => BU12545_A0,
         A1 => BU12545_A1,
         A2 => BU12545_A2,
         A3 => BU12545_A3,
         Q => BU12545_Q
      );

   BU12546_D <= n78;
   BU12546_CE <= n6861;
   BU12546_CLK <= n183;
   BU12546_A0 <= n6857;
   BU12546_A1 <= n6858;
   BU12546_A2 <= n6859;
   BU12546_A3 <= n6860;
   n6742 <= BU12546_Q;
   BU12546 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12546_D,
         CE => BU12546_CE,
         CLK => BU12546_CLK,
         A0 => BU12546_A0,
         A1 => BU12546_A1,
         A2 => BU12546_A2,
         A3 => BU12546_A3,
         Q => BU12546_Q
      );

   BU12547_D <= n79;
   BU12547_CE <= n6861;
   BU12547_CLK <= n183;
   BU12547_A0 <= n6857;
   BU12547_A1 <= n6858;
   BU12547_A2 <= n6859;
   BU12547_A3 <= n6860;
   n6743 <= BU12547_Q;
   BU12547 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12547_D,
         CE => BU12547_CE,
         CLK => BU12547_CLK,
         A0 => BU12547_A0,
         A1 => BU12547_A1,
         A2 => BU12547_A2,
         A3 => BU12547_A3,
         Q => BU12547_Q
      );

   BU12548_D <= n80;
   BU12548_CE <= n6861;
   BU12548_CLK <= n183;
   BU12548_A0 <= n6857;
   BU12548_A1 <= n6858;
   BU12548_A2 <= n6859;
   BU12548_A3 <= n6860;
   n6744 <= BU12548_Q;
   BU12548 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12548_D,
         CE => BU12548_CE,
         CLK => BU12548_CLK,
         A0 => BU12548_A0,
         A1 => BU12548_A1,
         A2 => BU12548_A2,
         A3 => BU12548_A3,
         Q => BU12548_Q
      );

   BU12549_D <= n81;
   BU12549_CE <= n6861;
   BU12549_CLK <= n183;
   BU12549_A0 <= n6857;
   BU12549_A1 <= n6858;
   BU12549_A2 <= n6859;
   BU12549_A3 <= n6860;
   n6745 <= BU12549_Q;
   BU12549 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU12549_D,
         CE => BU12549_CE,
         CLK => BU12549_CLK,
         A0 => BU12549_A0,
         A1 => BU12549_A1,
         A2 => BU12549_A2,
         A3 => BU12549_A3,
         Q => BU12549_Q
      );

   n6857 <= BU12550_Q(0);
   n6858 <= BU12550_Q(1);
   n6859 <= BU12550_Q(2);
   n6860 <= BU12550_Q(3);
   BU12550_CLK <= n183;
   BU12550_UP <= n6861;
   BU12550_CE <= n6862;
   BU12550 : C_COUNTER_BINARY_V5_0
      GENERIC MAP (
         c_count_mode => 2,
         c_has_aset => 0,
         c_load_enable => 0,
         c_load_low => 0,
         c_count_to => "0000",
         c_sync_priority => 0,
         c_has_iv => 0,
         c_has_sclr => 0,
         c_restrict_count => 0,
         c_width => 4,
         c_has_q_thresh1 => 0,
         c_enable_rlocs => 0,
         c_has_q_thresh0 => 0,
         c_thresh1_value => "0000",
         c_has_load => 0,
         c_has_up => 0,
         c_thresh_early => 0,
         c_has_thresh1 => 0,
         c_has_thresh0 => 0,
         c_ainit_val => "0000",
         c_has_ce => 1,
         c_pipe_stages => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0000",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_count_by => "0001",
         c_has_l => 0,
         c_thresh0_value => "0000"
      )
      PORT MAP (
         Q => BU12550_Q,
         CLK => BU12550_CLK,
         UP => BU12550_UP,
         CE => BU12550_CE
      );

   BU12579_I0 <= n6746;
   BU12579_I1 <= n6861;
   BU12579_I2 <= n6747;
   BU12579_I3 <= n6863;
   n6862 <= BU12579_O;
   BU12579 : LUT4
      GENERIC MAP (
         INIT  => X"4060"
      )
      PORT MAP (
         I0 => BU12579_I0,
         I1 => BU12579_I1,
         I2 => BU12579_I2,
         I3 => BU12579_I3,
         O => BU12579_O
      );

   BU12583_I0 <= n6747;
   BU12583_I1 <= n6863;
   BU12583_I2 <= n6861;
   BU12583_I3 <= n6746;
   n7206 <= BU12583_O;
   BU12583 : LUT4
      GENERIC MAP (
         INIT  => X"e2ea"
      )
      PORT MAP (
         I0 => BU12583_I0,
         I1 => BU12583_I1,
         I2 => BU12583_I2,
         I3 => BU12583_I3,
         O => BU12583_O
      );

   BU12584_D <= n7206;
   BU12584_C <= n183;
   BU12584_CE <= '1';
   n6747 <= BU12584_Q;
   BU12584 : FDE
      PORT MAP (
         D => BU12584_D,
         C => BU12584_C,
         CE => BU12584_CE,
         Q => BU12584_Q
      );

   BU12587_I0 <= n6857;
   BU12587_I1 <= n6858;
   BU12587_I2 <= n6859;
   BU12587_I3 <= n6860;
   n6863 <= BU12587_O;
   BU12587 : LUT4
      GENERIC MAP (
         INIT  => X"0001"
      )
      PORT MAP (
         I0 => BU12587_I0,
         I1 => BU12587_I1,
         I2 => BU12587_I2,
         I3 => BU12587_I3,
         O => BU12587_O
      );

   BU12588_ND <= n6747;
   n6791 <= BU12588_RDY;
   BU12588_CLK <= n183;
   n6719 <= BU12588_RFD;
   BU12588_DIN(0) <= n6720;
   BU12588_DIN(1) <= n6721;
   BU12588_DIN(2) <= n6722;
   BU12588_DIN(3) <= n6723;
   BU12588_DIN(4) <= n6724;
   BU12588_DIN(5) <= n6725;
   BU12588_DIN(6) <= n6726;
   BU12588_DIN(7) <= n6727;
   BU12588_DIN(8) <= n6728;
   BU12588_DIN(9) <= n6729;
   BU12588_DIN(10) <= n6730;
   BU12588_DIN(11) <= n6731;
   BU12588_DIN(12) <= n6732;
   BU12588_DIN(13) <= n6733;
   BU12588_DIN(14) <= n6734;
   BU12588_DIN(15) <= n6735;
   BU12588_DIN(16) <= n6736;
   BU12588_DIN(17) <= n6737;
   BU12588_DIN(18) <= n6738;
   BU12588_DIN(19) <= n6739;
   BU12588_DIN(20) <= n6740;
   BU12588_DIN(21) <= n6741;
   BU12588_DIN(22) <= n6742;
   BU12588_DIN(23) <= n6743;
   BU12588_DIN(24) <= n6744;
   BU12588_DIN(25) <= n6745;
   n6748 <= BU12588_DOUT(0);
   n6749 <= BU12588_DOUT(1);
   n6750 <= BU12588_DOUT(2);
   n6751 <= BU12588_DOUT(3);
   n6752 <= BU12588_DOUT(4);
   n6753 <= BU12588_DOUT(5);
   n6754 <= BU12588_DOUT(6);
   n6755 <= BU12588_DOUT(7);
   n6756 <= BU12588_DOUT(8);
   n6757 <= BU12588_DOUT(9);
   n6758 <= BU12588_DOUT(10);
   n6759 <= BU12588_DOUT(11);
   n6760 <= BU12588_DOUT(12);
   n6761 <= BU12588_DOUT(13);
   n6762 <= BU12588_DOUT(14);
   n6763 <= BU12588_DOUT(15);
   n6764 <= BU12588_DOUT(16);
   n6765 <= BU12588_DOUT(17);
   n6766 <= BU12588_DOUT(18);
   n6767 <= BU12588_DOUT(19);
   n6768 <= BU12588_DOUT(20);
   n6769 <= BU12588_DOUT(21);
   n6770 <= BU12588_DOUT(22);
   n6771 <= BU12588_DOUT(23);
   n6772 <= BU12588_DOUT(24);
   n6773 <= BU12588_DOUT(25);
   n6774 <= BU12588_DOUT(26);
   n6775 <= BU12588_DOUT(27);
   n6776 <= BU12588_DOUT(28);
   n6777 <= BU12588_DOUT(29);
   n6778 <= BU12588_DOUT(30);
   n6779 <= BU12588_DOUT(31);
   n6780 <= BU12588_DOUT(32);
   n6781 <= BU12588_DOUT(33);
   n6782 <= BU12588_DOUT(34);
   n6783 <= BU12588_DOUT(35);
   n6784 <= BU12588_DOUT(36);
   n6785 <= BU12588_DOUT(37);
   n6786 <= BU12588_DOUT(38);
   n6787 <= BU12588_DOUT(39);
   n6788 <= BU12588_DOUT(40);
   n6789 <= BU12588_DOUT(41);
   n6790 <= BU12588_DOUT(42);
   BU12588 : C_DA_FIR_V7_0
      GENERIC MAP (
         c_has_sout_r => 0,
         c_result_width => 43,
         c_reload_delay => 401,
         c_data_type => 0,
         c_filter_type => 0,
         c_channels => 2,
         c_response => 0,
         c_has_sout_f => 0,
         c_reg_output => 0,
         c_taps => 45,
         c_data_width => 26,
         c_enable_rlocs => 0,
         c_coeff_type => 0,
         c_reload_mem_type => 2,
         c_has_sin_r => 0,
         c_reload => 0,
         c_baat => 6,
         c_latency => 15,
         c_coeff_width => 16,
         c_optimize => 1,
         c_use_model_func => 0,
         c_zpf => 1,
         c_has_sin_f => 0,
         c_shape => 0,
         c_saturate => 0,
         c_has_sel_o => 0,
         c_mem_init_file => "myddc_CFIR.mif",
         c_polyphase_factor => 1,
         c_has_sel_i => 0,
         c_has_reset => 0
      )
      PORT MAP (
         ND => BU12588_ND,
         RDY => BU12588_RDY,
         CLK => BU12588_CLK,
         RFD => BU12588_RFD,
         DIN => BU12588_DIN,
         DOUT => BU12588_DOUT
      );

   BU19118_I(0) <= n6748;
   BU19118_I(1) <= n6749;
   BU19118_I(2) <= n6750;
   BU19118_I(3) <= n6751;
   BU19118_I(4) <= n6752;
   BU19118_I(5) <= n6753;
   BU19118_I(6) <= n6754;
   BU19118_I(7) <= n6755;
   BU19118_I(8) <= n6756;
   BU19118_I(9) <= n6757;
   BU19118_I(10) <= n6758;
   BU19118_I(11) <= n6759;
   BU19118_I(12) <= n6760;
   n7367 <= BU19118_O;
   BU19118 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 13,
         c_input_inv_mask => "0111111111111"
      )
      PORT MAP (
         I => BU19118_I,
         O => BU19118_O
      );

   BU19133_I0 <= n6761;
   BU19133_I1 <= n6760;
   BU19133_I2 <= n7367;
   BU19133_I3 <= '0';
   n7364 <= BU19133_O;
   BU19133 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU19133_I0,
         I1 => BU19133_I1,
         I2 => BU19133_I2,
         I3 => BU19133_I3,
         O => BU19133_O
      );

   BU19134_A(0) <= n6761;
   BU19134_A(1) <= n6762;
   BU19134_A(2) <= n6763;
   BU19134_A(3) <= n6764;
   BU19134_A(4) <= n6765;
   BU19134_A(5) <= n6766;
   BU19134_A(6) <= n6767;
   BU19134_A(7) <= n6768;
   BU19134_A(8) <= n6769;
   BU19134_A(9) <= n6770;
   BU19134_A(10) <= n6771;
   BU19134_A(11) <= n6772;
   BU19134_A(12) <= n6773;
   BU19134_A(13) <= n6774;
   BU19134_A(14) <= n6775;
   BU19134_A(15) <= n6776;
   BU19134_A(16) <= n6777;
   BU19134_A(17) <= n6778;
   BU19134_A(18) <= n6779;
   BU19134_A(19) <= n6780;
   BU19134_A(20) <= n6781;
   BU19134_A(21) <= n6782;
   BU19134_A(22) <= n6783;
   BU19134_A(23) <= n6784;
   BU19134_A(24) <= n6785;
   BU19134_A(25) <= n6786;
   BU19134_A(26) <= n6787;
   BU19134_A(27) <= n6788;
   BU19134_A(28) <= n6789;
   BU19134_A(29) <= n6790;
   BU19134_B(0) <= n7364;
   n7333 <= BU19134_S(0);
   n7334 <= BU19134_S(1);
   n7335 <= BU19134_S(2);
   n7336 <= BU19134_S(3);
   n7337 <= BU19134_S(4);
   n7338 <= BU19134_S(5);
   n7339 <= BU19134_S(6);
   n7340 <= BU19134_S(7);
   n7341 <= BU19134_S(8);
   n7342 <= BU19134_S(9);
   n7343 <= BU19134_S(10);
   n7344 <= BU19134_S(11);
   n7345 <= BU19134_S(12);
   n7346 <= BU19134_S(13);
   n7347 <= BU19134_S(14);
   n7348 <= BU19134_S(15);
   n7349 <= BU19134_S(16);
   n7350 <= BU19134_S(17);
   n7351 <= BU19134_S(18);
   n7352 <= BU19134_S(19);
   n7353 <= BU19134_S(20);
   n7354 <= BU19134_S(21);
   n7355 <= BU19134_S(22);
   n7356 <= BU19134_S(23);
   n7357 <= BU19134_S(24);
   n7358 <= BU19134_S(25);
   n7359 <= BU19134_S(26);
   n7360 <= BU19134_S(27);
   n7361 <= BU19134_S(28);
   n7362 <= BU19134_S(29);
   BU19134 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 30,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 31,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 30,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU19134_A,
         B => BU19134_B,
         S => BU19134_S
      );

   BU19259_I0 <= n6790;
   BU19259_I1 <= n6789;
   BU19259_I2 <= n7362;
   BU19259_I3 <= '0';
   n7381 <= BU19259_O;
   BU19259 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU19259_I0,
         I1 => BU19259_I1,
         I2 => BU19259_I2,
         I3 => BU19259_I3,
         O => BU19259_O
      );

   BU19261_I0 <= n6790;
   BU19261_I1 <= n7362;
   BU19261_I2 <= '0';
   BU19261_I3 <= '0';
   n7383 <= BU19261_O;
   BU19261 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU19261_I0,
         I1 => BU19261_I1,
         I2 => BU19261_I2,
         I3 => BU19261_I3,
         O => BU19261_O
      );

   BU19262_D(0) <= n7333;
   BU19262_D(1) <= n7334;
   BU19262_D(2) <= n7335;
   BU19262_D(3) <= n7336;
   BU19262_D(4) <= n7337;
   BU19262_D(5) <= n7338;
   BU19262_D(6) <= n7339;
   BU19262_D(7) <= n7340;
   BU19262_D(8) <= n7341;
   BU19262_D(9) <= n7342;
   BU19262_D(10) <= n7343;
   BU19262_D(11) <= n7344;
   BU19262_D(12) <= n7345;
   BU19262_D(13) <= n7346;
   BU19262_D(14) <= n7347;
   BU19262_D(15) <= n7348;
   BU19262_D(16) <= n7349;
   BU19262_D(17) <= n7350;
   BU19262_D(18) <= n7351;
   BU19262_D(19) <= n7352;
   BU19262_D(20) <= n7353;
   BU19262_D(21) <= n7354;
   BU19262_D(22) <= n7355;
   BU19262_D(23) <= n7356;
   BU19262_D(24) <= n7357;
   BU19262_D(25) <= n7358;
   BU19262_D(26) <= n7359;
   BU19262_D(27) <= n7360;
   BU19262_D(28) <= n7361;
   n82 <= BU19262_Q(0);
   n83 <= BU19262_Q(1);
   n84 <= BU19262_Q(2);
   n85 <= BU19262_Q(3);
   n86 <= BU19262_Q(4);
   n87 <= BU19262_Q(5);
   n88 <= BU19262_Q(6);
   n89 <= BU19262_Q(7);
   n90 <= BU19262_Q(8);
   n91 <= BU19262_Q(9);
   n92 <= BU19262_Q(10);
   n93 <= BU19262_Q(11);
   n94 <= BU19262_Q(12);
   n95 <= BU19262_Q(13);
   n96 <= BU19262_Q(14);
   n97 <= BU19262_Q(15);
   n98 <= BU19262_Q(16);
   n99 <= BU19262_Q(17);
   n100 <= BU19262_Q(18);
   n101 <= BU19262_Q(19);
   n102 <= BU19262_Q(20);
   n103 <= BU19262_Q(21);
   n104 <= BU19262_Q(22);
   n105 <= BU19262_Q(23);
   n106 <= BU19262_Q(24);
   n107 <= BU19262_Q(25);
   n108 <= BU19262_Q(26);
   n109 <= BU19262_Q(27);
   n110 <= BU19262_Q(28);
   BU19262_CLK <= n183;
   BU19262_SCLR <= n7381;
   BU19262_SSET <= n7383;
   BU19262 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 29,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU19262_D,
         Q => BU19262_Q,
         CLK => BU19262_CLK,
         SCLR => BU19262_SCLR,
         SSET => BU19262_SSET
      );

   BU19379_D(0) <= n7362;
   n111 <= BU19379_Q(0);
   BU19379_CLK <= n183;
   BU19379_SCLR <= n7383;
   BU19379_SSET <= n7381;
   BU19379 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU19379_D,
         Q => BU19379_Q,
         CLK => BU19379_CLK,
         SCLR => BU19379_SCLR,
         SSET => BU19379_SSET
      );

   BU19386_D <= n6791;
   BU19386_C <= n183;
   BU19386_CE <= '1';
   n112 <= BU19386_Q;
   BU19386 : FDE
      PORT MAP (
         D => BU19386_D,
         C => BU19386_C,
         CE => BU19386_CE,
         Q => BU19386_Q
      );

   BU19389_ND <= n112;
   n162 <= BU19389_RDY;
   BU19389_CLK <= n183;
   BU19389_DIN(0) <= n82;
   BU19389_DIN(1) <= n83;
   BU19389_DIN(2) <= n84;
   BU19389_DIN(3) <= n85;
   BU19389_DIN(4) <= n86;
   BU19389_DIN(5) <= n87;
   BU19389_DIN(6) <= n88;
   BU19389_DIN(7) <= n89;
   BU19389_DIN(8) <= n90;
   BU19389_DIN(9) <= n91;
   BU19389_DIN(10) <= n92;
   BU19389_DIN(11) <= n93;
   BU19389_DIN(12) <= n94;
   BU19389_DIN(13) <= n95;
   BU19389_DIN(14) <= n96;
   BU19389_DIN(15) <= n97;
   BU19389_DIN(16) <= n98;
   BU19389_DIN(17) <= n99;
   BU19389_DIN(18) <= n100;
   BU19389_DIN(19) <= n101;
   BU19389_DIN(20) <= n102;
   BU19389_DIN(21) <= n103;
   BU19389_DIN(22) <= n104;
   BU19389_DIN(23) <= n105;
   BU19389_DIN(24) <= n106;
   BU19389_DIN(25) <= n107;
   BU19389_DIN(26) <= n108;
   BU19389_DIN(27) <= n109;
   BU19389_DIN(28) <= n110;
   BU19389_DIN(29) <= n111;
   n163 <= BU19389_SEL_O(0);
   n113 <= BU19389_DOUT(0);
   n114 <= BU19389_DOUT(1);
   n115 <= BU19389_DOUT(2);
   n116 <= BU19389_DOUT(3);
   n117 <= BU19389_DOUT(4);
   n118 <= BU19389_DOUT(5);
   n119 <= BU19389_DOUT(6);
   n120 <= BU19389_DOUT(7);
   n121 <= BU19389_DOUT(8);
   n122 <= BU19389_DOUT(9);
   n123 <= BU19389_DOUT(10);
   n124 <= BU19389_DOUT(11);
   n125 <= BU19389_DOUT(12);
   n126 <= BU19389_DOUT(13);
   n127 <= BU19389_DOUT(14);
   n128 <= BU19389_DOUT(15);
   n129 <= BU19389_DOUT(16);
   n130 <= BU19389_DOUT(17);
   n131 <= BU19389_DOUT(18);
   n132 <= BU19389_DOUT(19);
   n133 <= BU19389_DOUT(20);
   n134 <= BU19389_DOUT(21);
   n135 <= BU19389_DOUT(22);
   n136 <= BU19389_DOUT(23);
   n137 <= BU19389_DOUT(24);
   n138 <= BU19389_DOUT(25);
   n139 <= BU19389_DOUT(26);
   n140 <= BU19389_DOUT(27);
   n141 <= BU19389_DOUT(28);
   n142 <= BU19389_DOUT(29);
   n143 <= BU19389_DOUT(30);
   n144 <= BU19389_DOUT(31);
   n145 <= BU19389_DOUT(32);
   n146 <= BU19389_DOUT(33);
   n147 <= BU19389_DOUT(34);
   n148 <= BU19389_DOUT(35);
   n149 <= BU19389_DOUT(36);
   n150 <= BU19389_DOUT(37);
   n151 <= BU19389_DOUT(38);
   n152 <= BU19389_DOUT(39);
   n153 <= BU19389_DOUT(40);
   n154 <= BU19389_DOUT(41);
   n155 <= BU19389_DOUT(42);
   n156 <= BU19389_DOUT(43);
   n157 <= BU19389_DOUT(44);
   n158 <= BU19389_DOUT(45);
   n159 <= BU19389_DOUT(46);
   n160 <= BU19389_DOUT(47);
   n161 <= BU19389_DOUT(48);
   BU19389 : C_DA_FIR_V7_0
      GENERIC MAP (
         c_has_sout_r => 0,
         c_result_width => 49,
         c_reload_delay => 657,
         c_data_type => 0,
         c_filter_type => 2,
         c_channels => 2,
         c_response => 0,
         c_has_sout_f => 0,
         c_reg_output => 0,
         c_taps => 55,
         c_data_width => 30,
         c_enable_rlocs => 0,
         c_coeff_type => 0,
         c_reload_mem_type => 2,
         c_has_sin_r => 0,
         c_reload => 0,
         c_baat => 2,
         c_latency => 26,
         c_coeff_width => 16,
         c_optimize => 1,
         c_use_model_func => 0,
         c_zpf => 1,
         c_has_sin_f => 0,
         c_shape => 0,
         c_saturate => 0,
         c_has_sel_o => 1,
         c_mem_init_file => "myddc_PFIR.mif",
         c_polyphase_factor => 5,
         c_has_sel_i => 0,
         c_has_reset => 0
      )
      PORT MAP (
         ND => BU19389_ND,
         RDY => BU19389_RDY,
         CLK => BU19389_CLK,
         RFD => BU19389_RFD,
         DIN => BU19389_DIN,
         SEL_O => BU19389_SEL_O,
         DOUT => BU19389_DOUT
      );

   BU25395_I0 <= n162;
   BU25395_I1 <= n163;
   BU25395_I2 <= '0';
   BU25395_I3 <= '0';
   n164 <= BU25395_O;
   BU25395 : LUT4
      GENERIC MAP (
         INIT  => X"2222"
      )
      PORT MAP (
         I0 => BU25395_I0,
         I1 => BU25395_I1,
         I2 => BU25395_I2,
         I3 => BU25395_I3,
         O => BU25395_O
      );

   BU25397_I0 <= n162;
   BU25397_I1 <= n163;
   BU25397_I2 <= '0';
   BU25397_I3 <= '0';
   n165 <= BU25397_O;
   BU25397 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU25397_I0,
         I1 => BU25397_I1,
         I2 => BU25397_I2,
         I3 => BU25397_I3,
         O => BU25397_O
      );

   BU25400_D <= n165;
   BU25400_C <= n183;
   BU25400_CE <= '1';
   n181 <= BU25400_Q;
   BU25400 : FDE
      PORT MAP (
         D => BU25400_D,
         C => BU25400_C,
         CE => BU25400_CE,
         Q => BU25400_Q
      );

   BU25405_I(0) <= n113;
   BU25405_I(1) <= n114;
   BU25405_I(2) <= n115;
   BU25405_I(3) <= n116;
   BU25405_I(4) <= n117;
   BU25405_I(5) <= n118;
   BU25405_I(6) <= n119;
   BU25405_I(7) <= n120;
   BU25405_I(8) <= n121;
   BU25405_I(9) <= n122;
   BU25405_I(10) <= n123;
   BU25405_I(11) <= n124;
   BU25405_I(12) <= n125;
   BU25405_I(13) <= n126;
   BU25405_I(14) <= n127;
   BU25405_I(15) <= n128;
   BU25405_I(16) <= n129;
   BU25405_I(17) <= n130;
   BU25405_I(18) <= n131;
   n8133 <= BU25405_O;
   BU25405 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 19,
         c_input_inv_mask => "0111111111111111111"
      )
      PORT MAP (
         I => BU25405_I,
         O => BU25405_O
      );

   BU25427_I0 <= n132;
   BU25427_I1 <= n131;
   BU25427_I2 <= n8133;
   BU25427_I3 <= '0';
   n8130 <= BU25427_O;
   BU25427 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU25427_I0,
         I1 => BU25427_I1,
         I2 => BU25427_I2,
         I3 => BU25427_I3,
         O => BU25427_O
      );

   BU25428_A(0) <= n132;
   BU25428_A(1) <= n133;
   BU25428_A(2) <= n134;
   BU25428_A(3) <= n135;
   BU25428_A(4) <= n136;
   BU25428_A(5) <= n137;
   BU25428_A(6) <= n138;
   BU25428_A(7) <= n139;
   BU25428_A(8) <= n140;
   BU25428_A(9) <= n141;
   BU25428_A(10) <= n142;
   BU25428_A(11) <= n143;
   BU25428_A(12) <= n144;
   BU25428_A(13) <= n145;
   BU25428_A(14) <= n146;
   BU25428_A(15) <= n147;
   BU25428_A(16) <= n148;
   BU25428_A(17) <= n149;
   BU25428_A(18) <= n150;
   BU25428_A(19) <= n151;
   BU25428_A(20) <= n152;
   BU25428_A(21) <= n153;
   BU25428_A(22) <= n154;
   BU25428_A(23) <= n155;
   BU25428_A(24) <= n156;
   BU25428_A(25) <= n157;
   BU25428_A(26) <= n158;
   BU25428_A(27) <= n159;
   BU25428_A(28) <= n160;
   BU25428_A(29) <= n161;
   BU25428_B(0) <= n8130;
   n8099 <= BU25428_S(0);
   n8100 <= BU25428_S(1);
   n8101 <= BU25428_S(2);
   n8102 <= BU25428_S(3);
   n8103 <= BU25428_S(4);
   n8104 <= BU25428_S(5);
   n8105 <= BU25428_S(6);
   n8106 <= BU25428_S(7);
   n8107 <= BU25428_S(8);
   n8108 <= BU25428_S(9);
   n8109 <= BU25428_S(10);
   n8110 <= BU25428_S(11);
   n8111 <= BU25428_S(12);
   n8112 <= BU25428_S(13);
   n8113 <= BU25428_S(14);
   n8114 <= BU25428_S(15);
   n8115 <= BU25428_S(16);
   n8116 <= BU25428_S(17);
   n8117 <= BU25428_S(18);
   n8118 <= BU25428_S(19);
   n8119 <= BU25428_S(20);
   n8120 <= BU25428_S(21);
   n8121 <= BU25428_S(22);
   n8122 <= BU25428_S(23);
   n8123 <= BU25428_S(24);
   n8124 <= BU25428_S(25);
   n8125 <= BU25428_S(26);
   n8126 <= BU25428_S(27);
   n8127 <= BU25428_S(28);
   n8128 <= BU25428_S(29);
   BU25428 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 30,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 31,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 30,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU25428_A,
         B => BU25428_B,
         S => BU25428_S
      );

   BU25553_I0 <= n161;
   BU25553_I1 <= n160;
   BU25553_I2 <= n8128;
   BU25553_I3 <= n164;
   n8153 <= BU25553_O;
   BU25553 : LUT4
      GENERIC MAP (
         INIT  => X"0200"
      )
      PORT MAP (
         I0 => BU25553_I0,
         I1 => BU25553_I1,
         I2 => BU25553_I2,
         I3 => BU25553_I3,
         O => BU25553_O
      );

   BU25555_I0 <= n161;
   BU25555_I1 <= n8128;
   BU25555_I2 <= n164;
   BU25555_I3 <= '0';
   n8155 <= BU25555_O;
   BU25555 : LUT4
      GENERIC MAP (
         INIT  => X"4040"
      )
      PORT MAP (
         I0 => BU25555_I0,
         I1 => BU25555_I1,
         I2 => BU25555_I2,
         I3 => BU25555_I3,
         O => BU25555_O
      );

   BU25556_D(0) <= n8099;
   BU25556_D(1) <= n8100;
   BU25556_D(2) <= n8101;
   BU25556_D(3) <= n8102;
   BU25556_D(4) <= n8103;
   BU25556_D(5) <= n8104;
   BU25556_D(6) <= n8105;
   BU25556_D(7) <= n8106;
   BU25556_D(8) <= n8107;
   BU25556_D(9) <= n8108;
   BU25556_D(10) <= n8109;
   BU25556_D(11) <= n8110;
   BU25556_D(12) <= n8111;
   BU25556_D(13) <= n8112;
   BU25556_D(14) <= n8113;
   BU25556_D(15) <= n8114;
   BU25556_D(16) <= n8115;
   BU25556_D(17) <= n8116;
   BU25556_D(18) <= n8117;
   BU25556_D(19) <= n8118;
   BU25556_D(20) <= n8119;
   BU25556_D(21) <= n8120;
   BU25556_D(22) <= n8121;
   BU25556_D(23) <= n8122;
   BU25556_D(24) <= n8123;
   BU25556_D(25) <= n8124;
   BU25556_D(26) <= n8125;
   BU25556_D(27) <= n8126;
   BU25556_D(28) <= n8127;
   n223 <= BU25556_Q(0);
   n224 <= BU25556_Q(1);
   n225 <= BU25556_Q(2);
   n226 <= BU25556_Q(3);
   n227 <= BU25556_Q(4);
   n228 <= BU25556_Q(5);
   n229 <= BU25556_Q(6);
   n230 <= BU25556_Q(7);
   n231 <= BU25556_Q(8);
   n232 <= BU25556_Q(9);
   n233 <= BU25556_Q(10);
   n234 <= BU25556_Q(11);
   n235 <= BU25556_Q(12);
   n236 <= BU25556_Q(13);
   n237 <= BU25556_Q(14);
   n238 <= BU25556_Q(15);
   n239 <= BU25556_Q(16);
   n240 <= BU25556_Q(17);
   n241 <= BU25556_Q(18);
   n242 <= BU25556_Q(19);
   n243 <= BU25556_Q(20);
   n244 <= BU25556_Q(21);
   n245 <= BU25556_Q(22);
   n246 <= BU25556_Q(23);
   n247 <= BU25556_Q(24);
   n248 <= BU25556_Q(25);
   n249 <= BU25556_Q(26);
   n250 <= BU25556_Q(27);
   n251 <= BU25556_Q(28);
   BU25556_CLK <= n183;
   BU25556_CE <= n164;
   BU25556_SCLR <= n8153;
   BU25556_SSET <= n8155;
   BU25556 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 29,
         c_has_ce => 1,
         c_sinit_val => "00000000000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU25556_D,
         Q => BU25556_Q,
         CLK => BU25556_CLK,
         CE => BU25556_CE,
         SCLR => BU25556_SCLR,
         SSET => BU25556_SSET
      );

   BU25676_D(0) <= n8128;
   n252 <= BU25676_Q(0);
   BU25676_CLK <= n183;
   BU25676_CE <= n164;
   BU25676_SCLR <= n8155;
   BU25676_SSET <= n8153;
   BU25676 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 1,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU25676_D,
         Q => BU25676_Q,
         CLK => BU25676_CLK,
         CE => BU25676_CE,
         SCLR => BU25676_SCLR,
         SSET => BU25676_SSET
      );

   BU25688_I(0) <= n113;
   BU25688_I(1) <= n114;
   BU25688_I(2) <= n115;
   BU25688_I(3) <= n116;
   BU25688_I(4) <= n117;
   BU25688_I(5) <= n118;
   BU25688_I(6) <= n119;
   BU25688_I(7) <= n120;
   BU25688_I(8) <= n121;
   BU25688_I(9) <= n122;
   BU25688_I(10) <= n123;
   BU25688_I(11) <= n124;
   BU25688_I(12) <= n125;
   BU25688_I(13) <= n126;
   BU25688_I(14) <= n127;
   BU25688_I(15) <= n128;
   BU25688_I(16) <= n129;
   BU25688_I(17) <= n130;
   BU25688_I(18) <= n131;
   n8735 <= BU25688_O;
   BU25688 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 19,
         c_input_inv_mask => "0111111111111111111"
      )
      PORT MAP (
         I => BU25688_I,
         O => BU25688_O
      );

   BU25710_I0 <= n132;
   BU25710_I1 <= n131;
   BU25710_I2 <= n8735;
   BU25710_I3 <= '0';
   n8732 <= BU25710_O;
   BU25710 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU25710_I0,
         I1 => BU25710_I1,
         I2 => BU25710_I2,
         I3 => BU25710_I3,
         O => BU25710_O
      );

   BU25711_A(0) <= n132;
   BU25711_A(1) <= n133;
   BU25711_A(2) <= n134;
   BU25711_A(3) <= n135;
   BU25711_A(4) <= n136;
   BU25711_A(5) <= n137;
   BU25711_A(6) <= n138;
   BU25711_A(7) <= n139;
   BU25711_A(8) <= n140;
   BU25711_A(9) <= n141;
   BU25711_A(10) <= n142;
   BU25711_A(11) <= n143;
   BU25711_A(12) <= n144;
   BU25711_A(13) <= n145;
   BU25711_A(14) <= n146;
   BU25711_A(15) <= n147;
   BU25711_A(16) <= n148;
   BU25711_A(17) <= n149;
   BU25711_A(18) <= n150;
   BU25711_A(19) <= n151;
   BU25711_A(20) <= n152;
   BU25711_A(21) <= n153;
   BU25711_A(22) <= n154;
   BU25711_A(23) <= n155;
   BU25711_A(24) <= n156;
   BU25711_A(25) <= n157;
   BU25711_A(26) <= n158;
   BU25711_A(27) <= n159;
   BU25711_A(28) <= n160;
   BU25711_A(29) <= n161;
   BU25711_B(0) <= n8732;
   n8701 <= BU25711_S(0);
   n8702 <= BU25711_S(1);
   n8703 <= BU25711_S(2);
   n8704 <= BU25711_S(3);
   n8705 <= BU25711_S(4);
   n8706 <= BU25711_S(5);
   n8707 <= BU25711_S(6);
   n8708 <= BU25711_S(7);
   n8709 <= BU25711_S(8);
   n8710 <= BU25711_S(9);
   n8711 <= BU25711_S(10);
   n8712 <= BU25711_S(11);
   n8713 <= BU25711_S(12);
   n8714 <= BU25711_S(13);
   n8715 <= BU25711_S(14);
   n8716 <= BU25711_S(15);
   n8717 <= BU25711_S(16);
   n8718 <= BU25711_S(17);
   n8719 <= BU25711_S(18);
   n8720 <= BU25711_S(19);
   n8721 <= BU25711_S(20);
   n8722 <= BU25711_S(21);
   n8723 <= BU25711_S(22);
   n8724 <= BU25711_S(23);
   n8725 <= BU25711_S(24);
   n8726 <= BU25711_S(25);
   n8727 <= BU25711_S(26);
   n8728 <= BU25711_S(27);
   n8729 <= BU25711_S(28);
   n8730 <= BU25711_S(29);
   BU25711 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 30,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 31,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 30,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU25711_A,
         B => BU25711_B,
         S => BU25711_S
      );

   BU25836_I0 <= n161;
   BU25836_I1 <= n160;
   BU25836_I2 <= n8730;
   BU25836_I3 <= n165;
   n8755 <= BU25836_O;
   BU25836 : LUT4
      GENERIC MAP (
         INIT  => X"0200"
      )
      PORT MAP (
         I0 => BU25836_I0,
         I1 => BU25836_I1,
         I2 => BU25836_I2,
         I3 => BU25836_I3,
         O => BU25836_O
      );

   BU25838_I0 <= n161;
   BU25838_I1 <= n8730;
   BU25838_I2 <= n165;
   BU25838_I3 <= '0';
   n8757 <= BU25838_O;
   BU25838 : LUT4
      GENERIC MAP (
         INIT  => X"4040"
      )
      PORT MAP (
         I0 => BU25838_I0,
         I1 => BU25838_I1,
         I2 => BU25838_I2,
         I3 => BU25838_I3,
         O => BU25838_O
      );

   BU25839_D(0) <= n8701;
   BU25839_D(1) <= n8702;
   BU25839_D(2) <= n8703;
   BU25839_D(3) <= n8704;
   BU25839_D(4) <= n8705;
   BU25839_D(5) <= n8706;
   BU25839_D(6) <= n8707;
   BU25839_D(7) <= n8708;
   BU25839_D(8) <= n8709;
   BU25839_D(9) <= n8710;
   BU25839_D(10) <= n8711;
   BU25839_D(11) <= n8712;
   BU25839_D(12) <= n8713;
   BU25839_D(13) <= n8714;
   BU25839_D(14) <= n8715;
   BU25839_D(15) <= n8716;
   BU25839_D(16) <= n8717;
   BU25839_D(17) <= n8718;
   BU25839_D(18) <= n8719;
   BU25839_D(19) <= n8720;
   BU25839_D(20) <= n8721;
   BU25839_D(21) <= n8722;
   BU25839_D(22) <= n8723;
   BU25839_D(23) <= n8724;
   BU25839_D(24) <= n8725;
   BU25839_D(25) <= n8726;
   BU25839_D(26) <= n8727;
   BU25839_D(27) <= n8728;
   BU25839_D(28) <= n8729;
   n253 <= BU25839_Q(0);
   n254 <= BU25839_Q(1);
   n255 <= BU25839_Q(2);
   n256 <= BU25839_Q(3);
   n257 <= BU25839_Q(4);
   n258 <= BU25839_Q(5);
   n259 <= BU25839_Q(6);
   n260 <= BU25839_Q(7);
   n261 <= BU25839_Q(8);
   n262 <= BU25839_Q(9);
   n263 <= BU25839_Q(10);
   n264 <= BU25839_Q(11);
   n265 <= BU25839_Q(12);
   n266 <= BU25839_Q(13);
   n267 <= BU25839_Q(14);
   n268 <= BU25839_Q(15);
   n269 <= BU25839_Q(16);
   n270 <= BU25839_Q(17);
   n271 <= BU25839_Q(18);
   n272 <= BU25839_Q(19);
   n273 <= BU25839_Q(20);
   n274 <= BU25839_Q(21);
   n275 <= BU25839_Q(22);
   n276 <= BU25839_Q(23);
   n277 <= BU25839_Q(24);
   n278 <= BU25839_Q(25);
   n279 <= BU25839_Q(26);
   n280 <= BU25839_Q(27);
   n281 <= BU25839_Q(28);
   BU25839_CLK <= n183;
   BU25839_CE <= n165;
   BU25839_SCLR <= n8755;
   BU25839_SSET <= n8757;
   BU25839 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 29,
         c_has_ce => 1,
         c_sinit_val => "00000000000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU25839_D,
         Q => BU25839_Q,
         CLK => BU25839_CLK,
         CE => BU25839_CE,
         SCLR => BU25839_SCLR,
         SSET => BU25839_SSET
      );

   BU25959_D(0) <= n8730;
   n282 <= BU25959_Q(0);
   BU25959_CLK <= n183;
   BU25959_CE <= n165;
   BU25959_SCLR <= n8757;
   BU25959_SSET <= n8755;
   BU25959 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 1,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU25959_D,
         Q => BU25959_Q,
         CLK => BU25959_CLK,
         CE => BU25959_CE,
         SCLR => BU25959_SCLR,
         SSET => BU25959_SSET
      );


END xilinx;


-- synthesis translate_on
