--------------------------------------------------------------------------------
--     This file is owned and controlled by Xilinx and must be used           --
--     solely for design, simulation, implementation and creation of          --
--     design files limited to Xilinx devices or technologies. Use            --
--     with non-Xilinx devices or technologies is expressly prohibited        --
--     and immediately terminates your license.                               --
--                                                                            --
--     XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS"          --
--     SOLELY FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR                --
--     XILINX DEVICES.  BY PROVIDING THIS DESIGN, CODE, OR INFORMATION        --
--     AS ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE, APPLICATION            --
--     OR STANDARD, XILINX IS MAKING NO REPRESENTATION THAT THIS              --
--     IMPLEMENTATION IS FREE FROM ANY CLAIMS OF INFRINGEMENT,                --
--     AND YOU ARE RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY REQUIRE       --
--     FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY DISCLAIMS ANY               --
--     WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE                --
--     IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR         --
--     REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF        --
--     INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS        --
--     FOR A PARTICULAR PURPOSE.                                              --
--                                                                            --
--     Xilinx products are not intended for use in life support               --
--     appliances, devices, or systems. Use in such applications are          --
--     expressly prohibited.                                                  --
--                                                                            --
--     (c) Copyright 1995-2004 Xilinx, Inc.                                   --
--     All rights reserved.                                                   --
--------------------------------------------------------------------------------

-- synopsys translate_off
LIBRARY std, ieee;
USE std.standard.ALL;
USE ieee.std_logic_1164.ALL;

LIBRARY unisim;
USE unisim.vcomponents.ALL;


LIBRARY XilinxCoreLib;
USE XilinxCoreLib.c_addsub_v5_0_comp.ALL;
USE XilinxCoreLib.c_da_fir_v7_0_comp.ALL;
USE XilinxCoreLib.c_mux_bus_v5_0_comp.ALL;
USE XilinxCoreLib.c_cic_v3_0_comp.ALL;
USE XilinxCoreLib.c_reg_fd_v5_0_comp.ALL;
USE XilinxCoreLib.c_dds_v4_1_comp.ALL;
USE XilinxCoreLib.c_shift_ram_v5_0_comp.ALL;
USE XilinxCoreLib.mult_gen_v5_0_comp.ALL;
USE XilinxCoreLib.c_gate_bit_v5_0_comp.ALL;

ENTITY ddcv1_0 IS
   PORT (
      DIN : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
      ND : IN STD_LOGIC;
      CLK : IN STD_LOGIC;
      ADDR : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      LD_DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      WE : IN STD_LOGIC;
      SEL : IN STD_LOGIC;
      RDY : OUT STD_LOGIC;
      RFD : OUT STD_LOGIC;
      DOUT_I : OUT STD_LOGIC_VECTOR(29 DOWNTO 0);
      DOUT_Q : OUT STD_LOGIC_VECTOR(29 DOWNTO 0)   
);
END ddcv1_0;

ARCHITECTURE xilinx OF ddcv1_0 IS 

-- Signals for connecting to instantiations
   SIGNAL BU4_I0 : STD_LOGIC;
   SIGNAL BU4_I1 : STD_LOGIC;
   SIGNAL BU4_I2 : STD_LOGIC;
   SIGNAL BU4_I3 : STD_LOGIC;
   SIGNAL BU4_O : STD_LOGIC;
   SIGNAL BU8_I0 : STD_LOGIC;
   SIGNAL BU8_I1 : STD_LOGIC;
   SIGNAL BU8_I2 : STD_LOGIC;
   SIGNAL BU8_I3 : STD_LOGIC;
   SIGNAL BU8_O : STD_LOGIC;
   SIGNAL BU10_I0 : STD_LOGIC;
   SIGNAL BU10_I1 : STD_LOGIC;
   SIGNAL BU10_I2 : STD_LOGIC;
   SIGNAL BU10_I3 : STD_LOGIC;
   SIGNAL BU10_O : STD_LOGIC;
   SIGNAL BU1292_D : STD_LOGIC;
   SIGNAL BU1292_C : STD_LOGIC;
   SIGNAL BU1292_CE : STD_LOGIC;
   SIGNAL BU1292_Q : STD_LOGIC;
   SIGNAL BU14_D : STD_LOGIC;
   SIGNAL BU14_CE : STD_LOGIC;
   SIGNAL BU14_CLK : STD_LOGIC;
   SIGNAL BU14_A0 : STD_LOGIC;
   SIGNAL BU14_A1 : STD_LOGIC;
   SIGNAL BU14_A2 : STD_LOGIC;
   SIGNAL BU14_A3 : STD_LOGIC;
   SIGNAL BU14_Q : STD_LOGIC;
   SIGNAL BU16_D : STD_LOGIC;
   SIGNAL BU16_C : STD_LOGIC;
   SIGNAL BU16_CE : STD_LOGIC;
   SIGNAL BU16_Q : STD_LOGIC;
   SIGNAL BU17_D : STD_LOGIC;
   SIGNAL BU17_CE : STD_LOGIC;
   SIGNAL BU17_CLK : STD_LOGIC;
   SIGNAL BU17_A0 : STD_LOGIC;
   SIGNAL BU17_A1 : STD_LOGIC;
   SIGNAL BU17_A2 : STD_LOGIC;
   SIGNAL BU17_A3 : STD_LOGIC;
   SIGNAL BU17_Q : STD_LOGIC;
   SIGNAL BU19_D : STD_LOGIC;
   SIGNAL BU19_C : STD_LOGIC;
   SIGNAL BU19_CE : STD_LOGIC;
   SIGNAL BU19_Q : STD_LOGIC;
   SIGNAL BU20_D : STD_LOGIC;
   SIGNAL BU20_CE : STD_LOGIC;
   SIGNAL BU20_CLK : STD_LOGIC;
   SIGNAL BU20_A0 : STD_LOGIC;
   SIGNAL BU20_A1 : STD_LOGIC;
   SIGNAL BU20_A2 : STD_LOGIC;
   SIGNAL BU20_A3 : STD_LOGIC;
   SIGNAL BU20_Q : STD_LOGIC;
   SIGNAL BU22_D : STD_LOGIC;
   SIGNAL BU22_C : STD_LOGIC;
   SIGNAL BU22_CE : STD_LOGIC;
   SIGNAL BU22_Q : STD_LOGIC;
   SIGNAL BU23_D : STD_LOGIC;
   SIGNAL BU23_CE : STD_LOGIC;
   SIGNAL BU23_CLK : STD_LOGIC;
   SIGNAL BU23_A0 : STD_LOGIC;
   SIGNAL BU23_A1 : STD_LOGIC;
   SIGNAL BU23_A2 : STD_LOGIC;
   SIGNAL BU23_A3 : STD_LOGIC;
   SIGNAL BU23_Q : STD_LOGIC;
   SIGNAL BU25_D : STD_LOGIC;
   SIGNAL BU25_C : STD_LOGIC;
   SIGNAL BU25_CE : STD_LOGIC;
   SIGNAL BU25_Q : STD_LOGIC;
   SIGNAL BU26_D : STD_LOGIC;
   SIGNAL BU26_CE : STD_LOGIC;
   SIGNAL BU26_CLK : STD_LOGIC;
   SIGNAL BU26_A0 : STD_LOGIC;
   SIGNAL BU26_A1 : STD_LOGIC;
   SIGNAL BU26_A2 : STD_LOGIC;
   SIGNAL BU26_A3 : STD_LOGIC;
   SIGNAL BU26_Q : STD_LOGIC;
   SIGNAL BU28_D : STD_LOGIC;
   SIGNAL BU28_C : STD_LOGIC;
   SIGNAL BU28_CE : STD_LOGIC;
   SIGNAL BU28_Q : STD_LOGIC;
   SIGNAL BU29_D : STD_LOGIC;
   SIGNAL BU29_CE : STD_LOGIC;
   SIGNAL BU29_CLK : STD_LOGIC;
   SIGNAL BU29_A0 : STD_LOGIC;
   SIGNAL BU29_A1 : STD_LOGIC;
   SIGNAL BU29_A2 : STD_LOGIC;
   SIGNAL BU29_A3 : STD_LOGIC;
   SIGNAL BU29_Q : STD_LOGIC;
   SIGNAL BU31_D : STD_LOGIC;
   SIGNAL BU31_C : STD_LOGIC;
   SIGNAL BU31_CE : STD_LOGIC;
   SIGNAL BU31_Q : STD_LOGIC;
   SIGNAL BU32_D : STD_LOGIC;
   SIGNAL BU32_CE : STD_LOGIC;
   SIGNAL BU32_CLK : STD_LOGIC;
   SIGNAL BU32_A0 : STD_LOGIC;
   SIGNAL BU32_A1 : STD_LOGIC;
   SIGNAL BU32_A2 : STD_LOGIC;
   SIGNAL BU32_A3 : STD_LOGIC;
   SIGNAL BU32_Q : STD_LOGIC;
   SIGNAL BU34_D : STD_LOGIC;
   SIGNAL BU34_C : STD_LOGIC;
   SIGNAL BU34_CE : STD_LOGIC;
   SIGNAL BU34_Q : STD_LOGIC;
   SIGNAL BU35_D : STD_LOGIC;
   SIGNAL BU35_CE : STD_LOGIC;
   SIGNAL BU35_CLK : STD_LOGIC;
   SIGNAL BU35_A0 : STD_LOGIC;
   SIGNAL BU35_A1 : STD_LOGIC;
   SIGNAL BU35_A2 : STD_LOGIC;
   SIGNAL BU35_A3 : STD_LOGIC;
   SIGNAL BU35_Q : STD_LOGIC;
   SIGNAL BU37_D : STD_LOGIC;
   SIGNAL BU37_C : STD_LOGIC;
   SIGNAL BU37_CE : STD_LOGIC;
   SIGNAL BU37_Q : STD_LOGIC;
   SIGNAL BU38_D : STD_LOGIC;
   SIGNAL BU38_CE : STD_LOGIC;
   SIGNAL BU38_CLK : STD_LOGIC;
   SIGNAL BU38_A0 : STD_LOGIC;
   SIGNAL BU38_A1 : STD_LOGIC;
   SIGNAL BU38_A2 : STD_LOGIC;
   SIGNAL BU38_A3 : STD_LOGIC;
   SIGNAL BU38_Q : STD_LOGIC;
   SIGNAL BU40_D : STD_LOGIC;
   SIGNAL BU40_C : STD_LOGIC;
   SIGNAL BU40_CE : STD_LOGIC;
   SIGNAL BU40_Q : STD_LOGIC;
   SIGNAL BU41_D : STD_LOGIC;
   SIGNAL BU41_CE : STD_LOGIC;
   SIGNAL BU41_CLK : STD_LOGIC;
   SIGNAL BU41_A0 : STD_LOGIC;
   SIGNAL BU41_A1 : STD_LOGIC;
   SIGNAL BU41_A2 : STD_LOGIC;
   SIGNAL BU41_A3 : STD_LOGIC;
   SIGNAL BU41_Q : STD_LOGIC;
   SIGNAL BU43_D : STD_LOGIC;
   SIGNAL BU43_C : STD_LOGIC;
   SIGNAL BU43_CE : STD_LOGIC;
   SIGNAL BU43_Q : STD_LOGIC;
   SIGNAL BU44_D : STD_LOGIC;
   SIGNAL BU44_CE : STD_LOGIC;
   SIGNAL BU44_CLK : STD_LOGIC;
   SIGNAL BU44_A0 : STD_LOGIC;
   SIGNAL BU44_A1 : STD_LOGIC;
   SIGNAL BU44_A2 : STD_LOGIC;
   SIGNAL BU44_A3 : STD_LOGIC;
   SIGNAL BU44_Q : STD_LOGIC;
   SIGNAL BU46_D : STD_LOGIC;
   SIGNAL BU46_C : STD_LOGIC;
   SIGNAL BU46_CE : STD_LOGIC;
   SIGNAL BU46_Q : STD_LOGIC;
   SIGNAL BU47_D : STD_LOGIC;
   SIGNAL BU47_CE : STD_LOGIC;
   SIGNAL BU47_CLK : STD_LOGIC;
   SIGNAL BU47_A0 : STD_LOGIC;
   SIGNAL BU47_A1 : STD_LOGIC;
   SIGNAL BU47_A2 : STD_LOGIC;
   SIGNAL BU47_A3 : STD_LOGIC;
   SIGNAL BU47_Q : STD_LOGIC;
   SIGNAL BU49_D : STD_LOGIC;
   SIGNAL BU49_C : STD_LOGIC;
   SIGNAL BU49_CE : STD_LOGIC;
   SIGNAL BU49_Q : STD_LOGIC;
   SIGNAL BU50_D : STD_LOGIC;
   SIGNAL BU50_CE : STD_LOGIC;
   SIGNAL BU50_CLK : STD_LOGIC;
   SIGNAL BU50_A0 : STD_LOGIC;
   SIGNAL BU50_A1 : STD_LOGIC;
   SIGNAL BU50_A2 : STD_LOGIC;
   SIGNAL BU50_A3 : STD_LOGIC;
   SIGNAL BU50_Q : STD_LOGIC;
   SIGNAL BU52_D : STD_LOGIC;
   SIGNAL BU52_C : STD_LOGIC;
   SIGNAL BU52_CE : STD_LOGIC;
   SIGNAL BU52_Q : STD_LOGIC;
   SIGNAL BU53_D : STD_LOGIC;
   SIGNAL BU53_CE : STD_LOGIC;
   SIGNAL BU53_CLK : STD_LOGIC;
   SIGNAL BU53_A0 : STD_LOGIC;
   SIGNAL BU53_A1 : STD_LOGIC;
   SIGNAL BU53_A2 : STD_LOGIC;
   SIGNAL BU53_A3 : STD_LOGIC;
   SIGNAL BU53_Q : STD_LOGIC;
   SIGNAL BU55_D : STD_LOGIC;
   SIGNAL BU55_C : STD_LOGIC;
   SIGNAL BU55_CE : STD_LOGIC;
   SIGNAL BU55_Q : STD_LOGIC;
   SIGNAL BU57_DATA : STD_LOGIC_VECTOR(31 DOWNTO 0);
   SIGNAL BU57_WE : STD_LOGIC;
   SIGNAL BU57_CLK : STD_LOGIC;
   SIGNAL BU57_CE : STD_LOGIC;
   SIGNAL BU57_RDY : STD_LOGIC;
   SIGNAL BU57_SINE : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU57_COSINE : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1294_I0 : STD_LOGIC;
   SIGNAL BU1294_I1 : STD_LOGIC;
   SIGNAL BU1294_I2 : STD_LOGIC;
   SIGNAL BU1294_I3 : STD_LOGIC;
   SIGNAL BU1294_O : STD_LOGIC;
   SIGNAL BU1296_clk : STD_LOGIC;
   SIGNAL BU1296_a : STD_LOGIC_VECTOR(13 DOWNTO 0);
   SIGNAL BU1296_b : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1296_o : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1296_q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1296_a_signed : STD_LOGIC;
   SIGNAL BU1296_loadb : STD_LOGIC;
   SIGNAL BU1296_load_done : STD_LOGIC;
   SIGNAL BU1296_swapb : STD_LOGIC;
   SIGNAL BU1296_ce : STD_LOGIC;
   SIGNAL BU1296_aclr : STD_LOGIC;
   SIGNAL BU1296_sclr : STD_LOGIC;
   SIGNAL BU1296_rfd : STD_LOGIC;
   SIGNAL BU1296_nd : STD_LOGIC;
   SIGNAL BU1296_rdy : STD_LOGIC;
   SIGNAL BU1517_I : STD_LOGIC_VECTOR(4 DOWNTO 0);
   SIGNAL BU1517_O : STD_LOGIC;
   SIGNAL BU1526_I0 : STD_LOGIC;
   SIGNAL BU1526_I1 : STD_LOGIC;
   SIGNAL BU1526_I2 : STD_LOGIC;
   SIGNAL BU1526_I3 : STD_LOGIC;
   SIGNAL BU1526_O : STD_LOGIC;
   SIGNAL BU1527_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU1527_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1527_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU1628_I0 : STD_LOGIC;
   SIGNAL BU1628_I1 : STD_LOGIC;
   SIGNAL BU1628_I2 : STD_LOGIC;
   SIGNAL BU1628_I3 : STD_LOGIC;
   SIGNAL BU1628_O : STD_LOGIC;
   SIGNAL BU1630_I0 : STD_LOGIC;
   SIGNAL BU1630_I1 : STD_LOGIC;
   SIGNAL BU1630_I2 : STD_LOGIC;
   SIGNAL BU1630_I3 : STD_LOGIC;
   SIGNAL BU1630_O : STD_LOGIC;
   SIGNAL BU1631_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU1631_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU1631_CLK : STD_LOGIC;
   SIGNAL BU1631_SCLR : STD_LOGIC;
   SIGNAL BU1631_SSET : STD_LOGIC;
   SIGNAL BU1724_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1724_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1724_CLK : STD_LOGIC;
   SIGNAL BU1724_SCLR : STD_LOGIC;
   SIGNAL BU1724_SSET : STD_LOGIC;
   SIGNAL BU1729_CLK : STD_LOGIC;
   SIGNAL BU1729_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1729_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1734_clk : STD_LOGIC;
   SIGNAL BU1734_a : STD_LOGIC_VECTOR(13 DOWNTO 0);
   SIGNAL BU1734_b : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU1734_o : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1734_q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU1734_a_signed : STD_LOGIC;
   SIGNAL BU1734_loadb : STD_LOGIC;
   SIGNAL BU1734_load_done : STD_LOGIC;
   SIGNAL BU1734_swapb : STD_LOGIC;
   SIGNAL BU1734_ce : STD_LOGIC;
   SIGNAL BU1734_aclr : STD_LOGIC;
   SIGNAL BU1734_sclr : STD_LOGIC;
   SIGNAL BU1734_rfd : STD_LOGIC;
   SIGNAL BU1734_nd : STD_LOGIC;
   SIGNAL BU1734_rdy : STD_LOGIC;
   SIGNAL BU1955_I : STD_LOGIC_VECTOR(4 DOWNTO 0);
   SIGNAL BU1955_O : STD_LOGIC;
   SIGNAL BU1964_I0 : STD_LOGIC;
   SIGNAL BU1964_I1 : STD_LOGIC;
   SIGNAL BU1964_I2 : STD_LOGIC;
   SIGNAL BU1964_I3 : STD_LOGIC;
   SIGNAL BU1964_O : STD_LOGIC;
   SIGNAL BU1965_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU1965_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU1965_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU2066_I0 : STD_LOGIC;
   SIGNAL BU2066_I1 : STD_LOGIC;
   SIGNAL BU2066_I2 : STD_LOGIC;
   SIGNAL BU2066_I3 : STD_LOGIC;
   SIGNAL BU2066_O : STD_LOGIC;
   SIGNAL BU2068_I0 : STD_LOGIC;
   SIGNAL BU2068_I1 : STD_LOGIC;
   SIGNAL BU2068_I2 : STD_LOGIC;
   SIGNAL BU2068_I3 : STD_LOGIC;
   SIGNAL BU2068_O : STD_LOGIC;
   SIGNAL BU2069_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2069_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2069_CLK : STD_LOGIC;
   SIGNAL BU2069_SCLR : STD_LOGIC;
   SIGNAL BU2069_SSET : STD_LOGIC;
   SIGNAL BU2162_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2162_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2162_CLK : STD_LOGIC;
   SIGNAL BU2162_SCLR : STD_LOGIC;
   SIGNAL BU2162_SSET : STD_LOGIC;
   SIGNAL BU2457_D : STD_LOGIC;
   SIGNAL BU2457_C : STD_LOGIC;
   SIGNAL BU2457_CE : STD_LOGIC;
   SIGNAL BU2457_Q : STD_LOGIC;
   SIGNAL BU2461_I : STD_LOGIC_VECTOR(15 DOWNTO 0);
   SIGNAL BU2461_O : STD_LOGIC;
   SIGNAL BU2479_I0 : STD_LOGIC;
   SIGNAL BU2479_I1 : STD_LOGIC;
   SIGNAL BU2479_I2 : STD_LOGIC;
   SIGNAL BU2479_I3 : STD_LOGIC;
   SIGNAL BU2479_O : STD_LOGIC;
   SIGNAL BU2480_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2480_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2480_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU2581_I0 : STD_LOGIC;
   SIGNAL BU2581_I1 : STD_LOGIC;
   SIGNAL BU2581_I2 : STD_LOGIC;
   SIGNAL BU2581_I3 : STD_LOGIC;
   SIGNAL BU2581_O : STD_LOGIC;
   SIGNAL BU2583_I0 : STD_LOGIC;
   SIGNAL BU2583_I1 : STD_LOGIC;
   SIGNAL BU2583_I2 : STD_LOGIC;
   SIGNAL BU2583_I3 : STD_LOGIC;
   SIGNAL BU2583_O : STD_LOGIC;
   SIGNAL BU2584_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2584_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU2584_CLK : STD_LOGIC;
   SIGNAL BU2584_SCLR : STD_LOGIC;
   SIGNAL BU2584_SSET : STD_LOGIC;
   SIGNAL BU2677_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2677_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2677_CLK : STD_LOGIC;
   SIGNAL BU2677_SCLR : STD_LOGIC;
   SIGNAL BU2677_SSET : STD_LOGIC;
   SIGNAL BU6771_I : STD_LOGIC_VECTOR(15 DOWNTO 0);
   SIGNAL BU6771_O : STD_LOGIC;
   SIGNAL BU6789_I0 : STD_LOGIC;
   SIGNAL BU6789_I1 : STD_LOGIC;
   SIGNAL BU6789_I2 : STD_LOGIC;
   SIGNAL BU6789_I3 : STD_LOGIC;
   SIGNAL BU6789_O : STD_LOGIC;
   SIGNAL BU6790_A : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU6790_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU6790_S : STD_LOGIC_VECTOR(24 DOWNTO 0);
   SIGNAL BU6891_I0 : STD_LOGIC;
   SIGNAL BU6891_I1 : STD_LOGIC;
   SIGNAL BU6891_I2 : STD_LOGIC;
   SIGNAL BU6891_I3 : STD_LOGIC;
   SIGNAL BU6891_O : STD_LOGIC;
   SIGNAL BU6893_I0 : STD_LOGIC;
   SIGNAL BU6893_I1 : STD_LOGIC;
   SIGNAL BU6893_I2 : STD_LOGIC;
   SIGNAL BU6893_I3 : STD_LOGIC;
   SIGNAL BU6893_O : STD_LOGIC;
   SIGNAL BU6894_D : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU6894_Q : STD_LOGIC_VECTOR(22 DOWNTO 0);
   SIGNAL BU6894_CLK : STD_LOGIC;
   SIGNAL BU6894_SCLR : STD_LOGIC;
   SIGNAL BU6894_SSET : STD_LOGIC;
   SIGNAL BU6987_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU6987_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU6987_CLK : STD_LOGIC;
   SIGNAL BU6987_SCLR : STD_LOGIC;
   SIGNAL BU6987_SSET : STD_LOGIC;
   SIGNAL BU2173_D : STD_LOGIC;
   SIGNAL BU2173_C : STD_LOGIC;
   SIGNAL BU2173_CE : STD_LOGIC;
   SIGNAL BU2173_Q : STD_LOGIC;
   SIGNAL BU2175_D : STD_LOGIC;
   SIGNAL BU2175_C : STD_LOGIC;
   SIGNAL BU2175_CE : STD_LOGIC;
   SIGNAL BU2175_Q : STD_LOGIC;
   SIGNAL BU2177_D : STD_LOGIC;
   SIGNAL BU2177_C : STD_LOGIC;
   SIGNAL BU2177_CE : STD_LOGIC;
   SIGNAL BU2177_Q : STD_LOGIC;
   SIGNAL BU2179_D : STD_LOGIC;
   SIGNAL BU2179_C : STD_LOGIC;
   SIGNAL BU2179_CE : STD_LOGIC;
   SIGNAL BU2179_Q : STD_LOGIC;
   SIGNAL BU2181_D : STD_LOGIC;
   SIGNAL BU2181_C : STD_LOGIC;
   SIGNAL BU2181_CE : STD_LOGIC;
   SIGNAL BU2181_Q : STD_LOGIC;
   SIGNAL BU2183_D : STD_LOGIC;
   SIGNAL BU2183_C : STD_LOGIC;
   SIGNAL BU2183_CE : STD_LOGIC;
   SIGNAL BU2183_Q : STD_LOGIC;
   SIGNAL BU2185_D : STD_LOGIC;
   SIGNAL BU2185_C : STD_LOGIC;
   SIGNAL BU2185_CE : STD_LOGIC;
   SIGNAL BU2185_Q : STD_LOGIC;
   SIGNAL BU2187_D : STD_LOGIC;
   SIGNAL BU2187_C : STD_LOGIC;
   SIGNAL BU2187_CE : STD_LOGIC;
   SIGNAL BU2187_Q : STD_LOGIC;
   SIGNAL BU2189_D : STD_LOGIC;
   SIGNAL BU2189_C : STD_LOGIC;
   SIGNAL BU2189_CE : STD_LOGIC;
   SIGNAL BU2189_Q : STD_LOGIC;
   SIGNAL BU2191_D : STD_LOGIC;
   SIGNAL BU2191_C : STD_LOGIC;
   SIGNAL BU2191_CE : STD_LOGIC;
   SIGNAL BU2191_Q : STD_LOGIC;
   SIGNAL BU2193_D : STD_LOGIC;
   SIGNAL BU2193_C : STD_LOGIC;
   SIGNAL BU2193_CE : STD_LOGIC;
   SIGNAL BU2193_Q : STD_LOGIC;
   SIGNAL BU2195_D : STD_LOGIC;
   SIGNAL BU2195_C : STD_LOGIC;
   SIGNAL BU2195_CE : STD_LOGIC;
   SIGNAL BU2195_Q : STD_LOGIC;
   SIGNAL BU2197_D : STD_LOGIC;
   SIGNAL BU2197_C : STD_LOGIC;
   SIGNAL BU2197_CE : STD_LOGIC;
   SIGNAL BU2197_Q : STD_LOGIC;
   SIGNAL BU2199_D : STD_LOGIC;
   SIGNAL BU2199_C : STD_LOGIC;
   SIGNAL BU2199_CE : STD_LOGIC;
   SIGNAL BU2199_Q : STD_LOGIC;
   SIGNAL BU2201_D : STD_LOGIC;
   SIGNAL BU2201_C : STD_LOGIC;
   SIGNAL BU2201_CE : STD_LOGIC;
   SIGNAL BU2201_Q : STD_LOGIC;
   SIGNAL BU2203_D : STD_LOGIC;
   SIGNAL BU2203_C : STD_LOGIC;
   SIGNAL BU2203_CE : STD_LOGIC;
   SIGNAL BU2203_Q : STD_LOGIC;
   SIGNAL BU2205_D : STD_LOGIC;
   SIGNAL BU2205_C : STD_LOGIC;
   SIGNAL BU2205_CE : STD_LOGIC;
   SIGNAL BU2205_Q : STD_LOGIC;
   SIGNAL BU2207_D : STD_LOGIC;
   SIGNAL BU2207_C : STD_LOGIC;
   SIGNAL BU2207_CE : STD_LOGIC;
   SIGNAL BU2207_Q : STD_LOGIC;
   SIGNAL BU2209_D : STD_LOGIC;
   SIGNAL BU2209_C : STD_LOGIC;
   SIGNAL BU2209_CE : STD_LOGIC;
   SIGNAL BU2209_Q : STD_LOGIC;
   SIGNAL BU2211_D : STD_LOGIC;
   SIGNAL BU2211_C : STD_LOGIC;
   SIGNAL BU2211_CE : STD_LOGIC;
   SIGNAL BU2211_Q : STD_LOGIC;
   SIGNAL BU2213_D : STD_LOGIC;
   SIGNAL BU2213_C : STD_LOGIC;
   SIGNAL BU2213_CE : STD_LOGIC;
   SIGNAL BU2213_Q : STD_LOGIC;
   SIGNAL BU2215_D : STD_LOGIC;
   SIGNAL BU2215_C : STD_LOGIC;
   SIGNAL BU2215_CE : STD_LOGIC;
   SIGNAL BU2215_Q : STD_LOGIC;
   SIGNAL BU2217_D : STD_LOGIC;
   SIGNAL BU2217_C : STD_LOGIC;
   SIGNAL BU2217_CE : STD_LOGIC;
   SIGNAL BU2217_Q : STD_LOGIC;
   SIGNAL BU2219_D : STD_LOGIC;
   SIGNAL BU2219_C : STD_LOGIC;
   SIGNAL BU2219_CE : STD_LOGIC;
   SIGNAL BU2219_Q : STD_LOGIC;
   SIGNAL BU2220_MA : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_MB : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_S : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU2220_Q : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2220_CLK : STD_LOGIC;
   SIGNAL BU2448_D : STD_LOGIC;
   SIGNAL BU2448_C : STD_LOGIC;
   SIGNAL BU2448_CE : STD_LOGIC;
   SIGNAL BU2448_Q : STD_LOGIC;
   SIGNAL BU2452_I0 : STD_LOGIC;
   SIGNAL BU2452_I1 : STD_LOGIC;
   SIGNAL BU2452_I2 : STD_LOGIC;
   SIGNAL BU2452_I3 : STD_LOGIC;
   SIGNAL BU2452_O : STD_LOGIC;
   SIGNAL BU2453_D : STD_LOGIC;
   SIGNAL BU2453_C : STD_LOGIC;
   SIGNAL BU2453_CE : STD_LOGIC;
   SIGNAL BU2453_Q : STD_LOGIC;
   SIGNAL BU2682_DIN : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU2682_ND : STD_LOGIC;
   SIGNAL BU2682_RFD : STD_LOGIC;
   SIGNAL BU2682_CLK : STD_LOGIC;
   SIGNAL BU2682_DOUT : STD_LOGIC_VECTOR(39 DOWNTO 0);
   SIGNAL BU2682_RDY : STD_LOGIC;
   SIGNAL BU6992_DIN : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU6992_ND : STD_LOGIC;
   SIGNAL BU6992_RFD : STD_LOGIC;
   SIGNAL BU6992_CLK : STD_LOGIC;
   SIGNAL BU6992_DOUT : STD_LOGIC_VECTOR(39 DOWNTO 0);
   SIGNAL BU6992_RDY : STD_LOGIC;
   SIGNAL BU11080_ND : STD_LOGIC;
   SIGNAL BU11080_RDY : STD_LOGIC;
   SIGNAL BU11080_CLK : STD_LOGIC;
   SIGNAL BU11080_RFD : STD_LOGIC;
   SIGNAL BU11080_DIN : STD_LOGIC_VECTOR(23 DOWNTO 0);
   SIGNAL BU11080_DOUT : STD_LOGIC_VECTOR(41 DOWNTO 0);
   SIGNAL BU20456_I : STD_LOGIC_VECTOR(25 DOWNTO 0);
   SIGNAL BU20456_O : STD_LOGIC;
   SIGNAL BU20487_I0 : STD_LOGIC;
   SIGNAL BU20487_I1 : STD_LOGIC;
   SIGNAL BU20487_I2 : STD_LOGIC;
   SIGNAL BU20487_I3 : STD_LOGIC;
   SIGNAL BU20487_O : STD_LOGIC;
   SIGNAL BU20488_A : STD_LOGIC_VECTOR(15 DOWNTO 0);
   SIGNAL BU20488_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU20488_S : STD_LOGIC_VECTOR(16 DOWNTO 0);
   SIGNAL BU20557_I0 : STD_LOGIC;
   SIGNAL BU20557_I1 : STD_LOGIC;
   SIGNAL BU20557_I2 : STD_LOGIC;
   SIGNAL BU20557_I3 : STD_LOGIC;
   SIGNAL BU20557_O : STD_LOGIC;
   SIGNAL BU20559_I0 : STD_LOGIC;
   SIGNAL BU20559_I1 : STD_LOGIC;
   SIGNAL BU20559_I2 : STD_LOGIC;
   SIGNAL BU20559_I3 : STD_LOGIC;
   SIGNAL BU20559_O : STD_LOGIC;
   SIGNAL BU20560_D : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU20560_Q : STD_LOGIC_VECTOR(14 DOWNTO 0);
   SIGNAL BU20560_CLK : STD_LOGIC;
   SIGNAL BU20560_SCLR : STD_LOGIC;
   SIGNAL BU20560_SSET : STD_LOGIC;
   SIGNAL BU20621_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU20621_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU20621_CLK : STD_LOGIC;
   SIGNAL BU20621_SCLR : STD_LOGIC;
   SIGNAL BU20621_SSET : STD_LOGIC;
   SIGNAL BU20628_D : STD_LOGIC;
   SIGNAL BU20628_C : STD_LOGIC;
   SIGNAL BU20628_CE : STD_LOGIC;
   SIGNAL BU20628_Q : STD_LOGIC;
   SIGNAL BU20631_ND : STD_LOGIC;
   SIGNAL BU20631_RDY : STD_LOGIC;
   SIGNAL BU20631_CLK : STD_LOGIC;
   SIGNAL BU20631_RFD : STD_LOGIC;
   SIGNAL BU20631_DIN : STD_LOGIC_VECTOR(15 DOWNTO 0);
   SIGNAL BU20631_SEL_O : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU20631_DOUT : STD_LOGIC_VECTOR(33 DOWNTO 0);
   SIGNAL BU24197_I0 : STD_LOGIC;
   SIGNAL BU24197_I1 : STD_LOGIC;
   SIGNAL BU24197_I2 : STD_LOGIC;
   SIGNAL BU24197_I3 : STD_LOGIC;
   SIGNAL BU24197_O : STD_LOGIC;
   SIGNAL BU24199_I0 : STD_LOGIC;
   SIGNAL BU24199_I1 : STD_LOGIC;
   SIGNAL BU24199_I2 : STD_LOGIC;
   SIGNAL BU24199_I3 : STD_LOGIC;
   SIGNAL BU24199_O : STD_LOGIC;
   SIGNAL BU24202_D : STD_LOGIC;
   SIGNAL BU24202_C : STD_LOGIC;
   SIGNAL BU24202_CE : STD_LOGIC;
   SIGNAL BU24202_Q : STD_LOGIC;
   SIGNAL BU24207_I : STD_LOGIC_VECTOR(3 DOWNTO 0);
   SIGNAL BU24207_O : STD_LOGIC;
   SIGNAL BU24213_I0 : STD_LOGIC;
   SIGNAL BU24213_I1 : STD_LOGIC;
   SIGNAL BU24213_I2 : STD_LOGIC;
   SIGNAL BU24213_I3 : STD_LOGIC;
   SIGNAL BU24213_O : STD_LOGIC;
   SIGNAL BU24214_A : STD_LOGIC_VECTOR(29 DOWNTO 0);
   SIGNAL BU24214_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU24214_S : STD_LOGIC_VECTOR(30 DOWNTO 0);
   SIGNAL BU24339_I0 : STD_LOGIC;
   SIGNAL BU24339_I1 : STD_LOGIC;
   SIGNAL BU24339_I2 : STD_LOGIC;
   SIGNAL BU24339_I3 : STD_LOGIC;
   SIGNAL BU24339_O : STD_LOGIC;
   SIGNAL BU24341_I0 : STD_LOGIC;
   SIGNAL BU24341_I1 : STD_LOGIC;
   SIGNAL BU24341_I2 : STD_LOGIC;
   SIGNAL BU24341_I3 : STD_LOGIC;
   SIGNAL BU24341_O : STD_LOGIC;
   SIGNAL BU24342_D : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU24342_Q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU24342_CLK : STD_LOGIC;
   SIGNAL BU24342_CE : STD_LOGIC;
   SIGNAL BU24342_SCLR : STD_LOGIC;
   SIGNAL BU24342_SSET : STD_LOGIC;
   SIGNAL BU24462_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU24462_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU24462_CLK : STD_LOGIC;
   SIGNAL BU24462_CE : STD_LOGIC;
   SIGNAL BU24462_SCLR : STD_LOGIC;
   SIGNAL BU24462_SSET : STD_LOGIC;
   SIGNAL BU24474_I : STD_LOGIC_VECTOR(3 DOWNTO 0);
   SIGNAL BU24474_O : STD_LOGIC;
   SIGNAL BU24480_I0 : STD_LOGIC;
   SIGNAL BU24480_I1 : STD_LOGIC;
   SIGNAL BU24480_I2 : STD_LOGIC;
   SIGNAL BU24480_I3 : STD_LOGIC;
   SIGNAL BU24480_O : STD_LOGIC;
   SIGNAL BU24481_A : STD_LOGIC_VECTOR(29 DOWNTO 0);
   SIGNAL BU24481_B : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU24481_S : STD_LOGIC_VECTOR(30 DOWNTO 0);
   SIGNAL BU24606_I0 : STD_LOGIC;
   SIGNAL BU24606_I1 : STD_LOGIC;
   SIGNAL BU24606_I2 : STD_LOGIC;
   SIGNAL BU24606_I3 : STD_LOGIC;
   SIGNAL BU24606_O : STD_LOGIC;
   SIGNAL BU24608_I0 : STD_LOGIC;
   SIGNAL BU24608_I1 : STD_LOGIC;
   SIGNAL BU24608_I2 : STD_LOGIC;
   SIGNAL BU24608_I3 : STD_LOGIC;
   SIGNAL BU24608_O : STD_LOGIC;
   SIGNAL BU24609_D : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU24609_Q : STD_LOGIC_VECTOR(28 DOWNTO 0);
   SIGNAL BU24609_CLK : STD_LOGIC;
   SIGNAL BU24609_CE : STD_LOGIC;
   SIGNAL BU24609_SCLR : STD_LOGIC;
   SIGNAL BU24609_SSET : STD_LOGIC;
   SIGNAL BU24729_D : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU24729_Q : STD_LOGIC_VECTOR(0 DOWNTO 0);
   SIGNAL BU24729_CLK : STD_LOGIC;
   SIGNAL BU24729_CE : STD_LOGIC;
   SIGNAL BU24729_SCLR : STD_LOGIC;
   SIGNAL BU24729_SSET : STD_LOGIC;
   SIGNAL n0 : STD_LOGIC := '0';
   SIGNAL n1 : STD_LOGIC := '1';
   SIGNAL n2 : STD_LOGIC;
   SIGNAL n3 : STD_LOGIC;
   SIGNAL n4 : STD_LOGIC;
   SIGNAL n5 : STD_LOGIC;
   SIGNAL n6 : STD_LOGIC;
   SIGNAL n7 : STD_LOGIC;
   SIGNAL n8 : STD_LOGIC;
   SIGNAL n9 : STD_LOGIC;
   SIGNAL n10 : STD_LOGIC;
   SIGNAL n11 : STD_LOGIC;
   SIGNAL n12 : STD_LOGIC;
   SIGNAL n13 : STD_LOGIC;
   SIGNAL n14 : STD_LOGIC;
   SIGNAL n15 : STD_LOGIC;
   SIGNAL n16 : STD_LOGIC;
   SIGNAL n17 : STD_LOGIC;
   SIGNAL n18 : STD_LOGIC;
   SIGNAL n19 : STD_LOGIC;
   SIGNAL n20 : STD_LOGIC;
   SIGNAL n21 : STD_LOGIC;
   SIGNAL n22 : STD_LOGIC;
   SIGNAL n23 : STD_LOGIC;
   SIGNAL n24 : STD_LOGIC;
   SIGNAL n25 : STD_LOGIC;
   SIGNAL n26 : STD_LOGIC;
   SIGNAL n27 : STD_LOGIC;
   SIGNAL n28 : STD_LOGIC;
   SIGNAL n29 : STD_LOGIC;
   SIGNAL n30 : STD_LOGIC;
   SIGNAL n31 : STD_LOGIC;
   SIGNAL n32 : STD_LOGIC;
   SIGNAL n33 : STD_LOGIC;
   SIGNAL n34 : STD_LOGIC;
   SIGNAL n35 : STD_LOGIC;
   SIGNAL n36 : STD_LOGIC;
   SIGNAL n37 : STD_LOGIC;
   SIGNAL n38 : STD_LOGIC;
   SIGNAL n39 : STD_LOGIC;
   SIGNAL n40 : STD_LOGIC;
   SIGNAL n41 : STD_LOGIC;
   SIGNAL n42 : STD_LOGIC;
   SIGNAL n43 : STD_LOGIC;
   SIGNAL n44 : STD_LOGIC;
   SIGNAL n45 : STD_LOGIC;
   SIGNAL n46 : STD_LOGIC;
   SIGNAL n47 : STD_LOGIC;
   SIGNAL n48 : STD_LOGIC;
   SIGNAL n49 : STD_LOGIC;
   SIGNAL n50 : STD_LOGIC;
   SIGNAL n54 : STD_LOGIC;
   SIGNAL n55 : STD_LOGIC;
   SIGNAL n56 : STD_LOGIC;
   SIGNAL n57 : STD_LOGIC;
   SIGNAL n58 : STD_LOGIC;
   SIGNAL n59 : STD_LOGIC;
   SIGNAL n60 : STD_LOGIC;
   SIGNAL n61 : STD_LOGIC;
   SIGNAL n62 : STD_LOGIC;
   SIGNAL n63 : STD_LOGIC;
   SIGNAL n64 : STD_LOGIC;
   SIGNAL n65 : STD_LOGIC;
   SIGNAL n66 : STD_LOGIC;
   SIGNAL n67 : STD_LOGIC;
   SIGNAL n68 : STD_LOGIC;
   SIGNAL n69 : STD_LOGIC;
   SIGNAL n70 : STD_LOGIC;
   SIGNAL n71 : STD_LOGIC;
   SIGNAL n72 : STD_LOGIC;
   SIGNAL n73 : STD_LOGIC;
   SIGNAL n74 : STD_LOGIC;
   SIGNAL n75 : STD_LOGIC;
   SIGNAL n76 : STD_LOGIC;
   SIGNAL n77 : STD_LOGIC;
   SIGNAL n78 : STD_LOGIC;
   SIGNAL n79 : STD_LOGIC;
   SIGNAL n80 : STD_LOGIC;
   SIGNAL n81 : STD_LOGIC;
   SIGNAL n82 : STD_LOGIC;
   SIGNAL n83 : STD_LOGIC;
   SIGNAL n84 : STD_LOGIC;
   SIGNAL n85 : STD_LOGIC;
   SIGNAL n86 : STD_LOGIC;
   SIGNAL n87 : STD_LOGIC;
   SIGNAL n88 : STD_LOGIC;
   SIGNAL n89 : STD_LOGIC;
   SIGNAL n90 : STD_LOGIC;
   SIGNAL n91 : STD_LOGIC;
   SIGNAL n92 : STD_LOGIC;
   SIGNAL n93 : STD_LOGIC;
   SIGNAL n94 : STD_LOGIC;
   SIGNAL n95 : STD_LOGIC;
   SIGNAL n96 : STD_LOGIC;
   SIGNAL n97 : STD_LOGIC;
   SIGNAL n98 : STD_LOGIC;
   SIGNAL n99 : STD_LOGIC;
   SIGNAL n100 : STD_LOGIC;
   SIGNAL n101 : STD_LOGIC;
   SIGNAL n102 : STD_LOGIC;
   SIGNAL n103 : STD_LOGIC;
   SIGNAL n104 : STD_LOGIC;
   SIGNAL n105 : STD_LOGIC;
   SIGNAL n106 : STD_LOGIC;
   SIGNAL n107 : STD_LOGIC;
   SIGNAL n108 : STD_LOGIC;
   SIGNAL n109 : STD_LOGIC;
   SIGNAL n110 : STD_LOGIC;
   SIGNAL n111 : STD_LOGIC;
   SIGNAL n112 : STD_LOGIC;
   SIGNAL n113 : STD_LOGIC;
   SIGNAL n114 : STD_LOGIC;
   SIGNAL n115 : STD_LOGIC;
   SIGNAL n116 : STD_LOGIC;
   SIGNAL n117 : STD_LOGIC;
   SIGNAL n118 : STD_LOGIC;
   SIGNAL n119 : STD_LOGIC;
   SIGNAL n120 : STD_LOGIC;
   SIGNAL n121 : STD_LOGIC;
   SIGNAL n122 : STD_LOGIC;
   SIGNAL n123 : STD_LOGIC;
   SIGNAL n124 : STD_LOGIC;
   SIGNAL n125 : STD_LOGIC;
   SIGNAL n126 : STD_LOGIC;
   SIGNAL n127 : STD_LOGIC;
   SIGNAL n128 : STD_LOGIC;
   SIGNAL n129 : STD_LOGIC;
   SIGNAL n130 : STD_LOGIC;
   SIGNAL n131 : STD_LOGIC;
   SIGNAL n132 : STD_LOGIC;
   SIGNAL n133 : STD_LOGIC;
   SIGNAL n134 : STD_LOGIC;
   SIGNAL n135 : STD_LOGIC;
   SIGNAL n136 : STD_LOGIC;
   SIGNAL n137 : STD_LOGIC;
   SIGNAL n138 : STD_LOGIC;
   SIGNAL n139 : STD_LOGIC;
   SIGNAL n140 : STD_LOGIC;
   SIGNAL n141 : STD_LOGIC;
   SIGNAL n142 : STD_LOGIC;
   SIGNAL n143 : STD_LOGIC;
   SIGNAL n144 : STD_LOGIC;
   SIGNAL n145 : STD_LOGIC;
   SIGNAL n146 : STD_LOGIC;
   SIGNAL n147 : STD_LOGIC;
   SIGNAL n148 : STD_LOGIC;
   SIGNAL n149 : STD_LOGIC;
   SIGNAL n150 : STD_LOGIC;
   SIGNAL n151 : STD_LOGIC;
   SIGNAL n152 : STD_LOGIC;
   SIGNAL n153 : STD_LOGIC;
   SIGNAL n154 : STD_LOGIC;
   SIGNAL n155 : STD_LOGIC;
   SIGNAL n156 : STD_LOGIC;
   SIGNAL n157 : STD_LOGIC;
   SIGNAL n158 : STD_LOGIC;
   SIGNAL n159 : STD_LOGIC;
   SIGNAL n160 : STD_LOGIC;
   SIGNAL n161 : STD_LOGIC;
   SIGNAL n162 : STD_LOGIC;
   SIGNAL n163 : STD_LOGIC;
   SIGNAL n164 : STD_LOGIC;
   SIGNAL n165 : STD_LOGIC;
   SIGNAL n166 : STD_LOGIC;
   SIGNAL n167 : STD_LOGIC;
   SIGNAL n168 : STD_LOGIC;
   SIGNAL n169 : STD_LOGIC;
   SIGNAL n170 : STD_LOGIC;
   SIGNAL n171 : STD_LOGIC;
   SIGNAL n172 : STD_LOGIC;
   SIGNAL n173 : STD_LOGIC;
   SIGNAL n174 : STD_LOGIC;
   SIGNAL n175 : STD_LOGIC;
   SIGNAL n176 : STD_LOGIC;
   SIGNAL n177 : STD_LOGIC;
   SIGNAL n178 : STD_LOGIC;
   SIGNAL n179 : STD_LOGIC;
   SIGNAL n180 : STD_LOGIC;
   SIGNAL n181 : STD_LOGIC;
   SIGNAL n182 : STD_LOGIC;
   SIGNAL n183 : STD_LOGIC;
   SIGNAL n184 : STD_LOGIC;
   SIGNAL n185 : STD_LOGIC;
   SIGNAL n186 : STD_LOGIC;
   SIGNAL n187 : STD_LOGIC;
   SIGNAL n188 : STD_LOGIC;
   SIGNAL n189 : STD_LOGIC;
   SIGNAL n190 : STD_LOGIC;
   SIGNAL n191 : STD_LOGIC;
   SIGNAL n192 : STD_LOGIC;
   SIGNAL n193 : STD_LOGIC;
   SIGNAL n194 : STD_LOGIC;
   SIGNAL n195 : STD_LOGIC;
   SIGNAL n196 : STD_LOGIC;
   SIGNAL n197 : STD_LOGIC;
   SIGNAL n198 : STD_LOGIC;
   SIGNAL n199 : STD_LOGIC;
   SIGNAL n200 : STD_LOGIC;
   SIGNAL n201 : STD_LOGIC;
   SIGNAL n202 : STD_LOGIC;
   SIGNAL n203 : STD_LOGIC;
   SIGNAL n204 : STD_LOGIC;
   SIGNAL n205 : STD_LOGIC;
   SIGNAL n206 : STD_LOGIC;
   SIGNAL n207 : STD_LOGIC;
   SIGNAL n208 : STD_LOGIC;
   SIGNAL n209 : STD_LOGIC;
   SIGNAL n210 : STD_LOGIC;
   SIGNAL n211 : STD_LOGIC;
   SIGNAL n212 : STD_LOGIC;
   SIGNAL n213 : STD_LOGIC;
   SIGNAL n214 : STD_LOGIC;
   SIGNAL n215 : STD_LOGIC;
   SIGNAL n216 : STD_LOGIC;
   SIGNAL n217 : STD_LOGIC;
   SIGNAL n218 : STD_LOGIC;
   SIGNAL n219 : STD_LOGIC;
   SIGNAL n220 : STD_LOGIC;
   SIGNAL n221 : STD_LOGIC;
   SIGNAL n222 : STD_LOGIC;
   SIGNAL n223 : STD_LOGIC;
   SIGNAL n224 : STD_LOGIC;
   SIGNAL n225 : STD_LOGIC;
   SIGNAL n226 : STD_LOGIC;
   SIGNAL n227 : STD_LOGIC;
   SIGNAL n228 : STD_LOGIC;
   SIGNAL n229 : STD_LOGIC;
   SIGNAL n230 : STD_LOGIC;
   SIGNAL n231 : STD_LOGIC;
   SIGNAL n232 : STD_LOGIC;
   SIGNAL n233 : STD_LOGIC;
   SIGNAL n234 : STD_LOGIC;
   SIGNAL n235 : STD_LOGIC;
   SIGNAL n236 : STD_LOGIC;
   SIGNAL n237 : STD_LOGIC;
   SIGNAL n238 : STD_LOGIC;
   SIGNAL n239 : STD_LOGIC;
   SIGNAL n240 : STD_LOGIC;
   SIGNAL n241 : STD_LOGIC;
   SIGNAL n242 : STD_LOGIC;
   SIGNAL n243 : STD_LOGIC;
   SIGNAL n244 : STD_LOGIC;
   SIGNAL n245 : STD_LOGIC;
   SIGNAL n246 : STD_LOGIC;
   SIGNAL n247 : STD_LOGIC;
   SIGNAL n248 : STD_LOGIC;
   SIGNAL n249 : STD_LOGIC;
   SIGNAL n250 : STD_LOGIC;
   SIGNAL n251 : STD_LOGIC;
   SIGNAL n291 : STD_LOGIC;
   SIGNAL n338 : STD_LOGIC;
   SIGNAL n339 : STD_LOGIC;
   SIGNAL n340 : STD_LOGIC;
   SIGNAL n412 : STD_LOGIC;
   SIGNAL n413 : STD_LOGIC;
   SIGNAL n414 : STD_LOGIC;
   SIGNAL n415 : STD_LOGIC;
   SIGNAL n416 : STD_LOGIC;
   SIGNAL n417 : STD_LOGIC;
   SIGNAL n418 : STD_LOGIC;
   SIGNAL n419 : STD_LOGIC;
   SIGNAL n420 : STD_LOGIC;
   SIGNAL n421 : STD_LOGIC;
   SIGNAL n422 : STD_LOGIC;
   SIGNAL n423 : STD_LOGIC;
   SIGNAL n424 : STD_LOGIC;
   SIGNAL n425 : STD_LOGIC;
   SIGNAL n426 : STD_LOGIC;
   SIGNAL n457 : STD_LOGIC;
   SIGNAL n458 : STD_LOGIC;
   SIGNAL n459 : STD_LOGIC;
   SIGNAL n460 : STD_LOGIC;
   SIGNAL n461 : STD_LOGIC;
   SIGNAL n462 : STD_LOGIC;
   SIGNAL n463 : STD_LOGIC;
   SIGNAL n464 : STD_LOGIC;
   SIGNAL n465 : STD_LOGIC;
   SIGNAL n466 : STD_LOGIC;
   SIGNAL n467 : STD_LOGIC;
   SIGNAL n468 : STD_LOGIC;
   SIGNAL n469 : STD_LOGIC;
   SIGNAL n470 : STD_LOGIC;
   SIGNAL n471 : STD_LOGIC;
   SIGNAL n472 : STD_LOGIC;
   SIGNAL n473 : STD_LOGIC;
   SIGNAL n474 : STD_LOGIC;
   SIGNAL n475 : STD_LOGIC;
   SIGNAL n476 : STD_LOGIC;
   SIGNAL n477 : STD_LOGIC;
   SIGNAL n478 : STD_LOGIC;
   SIGNAL n479 : STD_LOGIC;
   SIGNAL n480 : STD_LOGIC;
   SIGNAL n481 : STD_LOGIC;
   SIGNAL n482 : STD_LOGIC;
   SIGNAL n483 : STD_LOGIC;
   SIGNAL n484 : STD_LOGIC;
   SIGNAL n485 : STD_LOGIC;
   SIGNAL n544 : STD_LOGIC;
   SIGNAL n574 : STD_LOGIC;
   SIGNAL n575 : STD_LOGIC;
   SIGNAL n576 : STD_LOGIC;
   SIGNAL n577 : STD_LOGIC;
   SIGNAL n578 : STD_LOGIC;
   SIGNAL n579 : STD_LOGIC;
   SIGNAL n580 : STD_LOGIC;
   SIGNAL n581 : STD_LOGIC;
   SIGNAL n582 : STD_LOGIC;
   SIGNAL n583 : STD_LOGIC;
   SIGNAL n584 : STD_LOGIC;
   SIGNAL n585 : STD_LOGIC;
   SIGNAL n586 : STD_LOGIC;
   SIGNAL n587 : STD_LOGIC;
   SIGNAL n616 : STD_LOGIC;
   SIGNAL n617 : STD_LOGIC;
   SIGNAL n618 : STD_LOGIC;
   SIGNAL n619 : STD_LOGIC;
   SIGNAL n620 : STD_LOGIC;
   SIGNAL n621 : STD_LOGIC;
   SIGNAL n622 : STD_LOGIC;
   SIGNAL n623 : STD_LOGIC;
   SIGNAL n624 : STD_LOGIC;
   SIGNAL n625 : STD_LOGIC;
   SIGNAL n626 : STD_LOGIC;
   SIGNAL n627 : STD_LOGIC;
   SIGNAL n628 : STD_LOGIC;
   SIGNAL n629 : STD_LOGIC;
   SIGNAL n630 : STD_LOGIC;
   SIGNAL n661 : STD_LOGIC;
   SIGNAL n662 : STD_LOGIC;
   SIGNAL n663 : STD_LOGIC;
   SIGNAL n664 : STD_LOGIC;
   SIGNAL n665 : STD_LOGIC;
   SIGNAL n666 : STD_LOGIC;
   SIGNAL n667 : STD_LOGIC;
   SIGNAL n668 : STD_LOGIC;
   SIGNAL n669 : STD_LOGIC;
   SIGNAL n670 : STD_LOGIC;
   SIGNAL n671 : STD_LOGIC;
   SIGNAL n672 : STD_LOGIC;
   SIGNAL n673 : STD_LOGIC;
   SIGNAL n674 : STD_LOGIC;
   SIGNAL n675 : STD_LOGIC;
   SIGNAL n676 : STD_LOGIC;
   SIGNAL n677 : STD_LOGIC;
   SIGNAL n678 : STD_LOGIC;
   SIGNAL n679 : STD_LOGIC;
   SIGNAL n680 : STD_LOGIC;
   SIGNAL n681 : STD_LOGIC;
   SIGNAL n682 : STD_LOGIC;
   SIGNAL n683 : STD_LOGIC;
   SIGNAL n684 : STD_LOGIC;
   SIGNAL n685 : STD_LOGIC;
   SIGNAL n686 : STD_LOGIC;
   SIGNAL n687 : STD_LOGIC;
   SIGNAL n688 : STD_LOGIC;
   SIGNAL n689 : STD_LOGIC;
   SIGNAL n924 : STD_LOGIC;
   SIGNAL n925 : STD_LOGIC;
   SIGNAL n926 : STD_LOGIC;
   SIGNAL n927 : STD_LOGIC;
   SIGNAL n928 : STD_LOGIC;
   SIGNAL n929 : STD_LOGIC;
   SIGNAL n930 : STD_LOGIC;
   SIGNAL n931 : STD_LOGIC;
   SIGNAL n932 : STD_LOGIC;
   SIGNAL n933 : STD_LOGIC;
   SIGNAL n934 : STD_LOGIC;
   SIGNAL n935 : STD_LOGIC;
   SIGNAL n936 : STD_LOGIC;
   SIGNAL n937 : STD_LOGIC;
   SIGNAL n1516 : STD_LOGIC;
   SIGNAL n1517 : STD_LOGIC;
   SIGNAL n1518 : STD_LOGIC;
   SIGNAL n1519 : STD_LOGIC;
   SIGNAL n1520 : STD_LOGIC;
   SIGNAL n1521 : STD_LOGIC;
   SIGNAL n1522 : STD_LOGIC;
   SIGNAL n1523 : STD_LOGIC;
   SIGNAL n1524 : STD_LOGIC;
   SIGNAL n1525 : STD_LOGIC;
   SIGNAL n1526 : STD_LOGIC;
   SIGNAL n1527 : STD_LOGIC;
   SIGNAL n1528 : STD_LOGIC;
   SIGNAL n1529 : STD_LOGIC;
   SIGNAL n1530 : STD_LOGIC;
   SIGNAL n1531 : STD_LOGIC;
   SIGNAL n1532 : STD_LOGIC;
   SIGNAL n1533 : STD_LOGIC;
   SIGNAL n1534 : STD_LOGIC;
   SIGNAL n1535 : STD_LOGIC;
   SIGNAL n1536 : STD_LOGIC;
   SIGNAL n1537 : STD_LOGIC;
   SIGNAL n1538 : STD_LOGIC;
   SIGNAL n1539 : STD_LOGIC;
   SIGNAL n1541 : STD_LOGIC;
   SIGNAL n1544 : STD_LOGIC;
   SIGNAL n1550 : STD_LOGIC;
   SIGNAL n1552 : STD_LOGIC;
   SIGNAL n2159 : STD_LOGIC;
   SIGNAL n2160 : STD_LOGIC;
   SIGNAL n2161 : STD_LOGIC;
   SIGNAL n2162 : STD_LOGIC;
   SIGNAL n2163 : STD_LOGIC;
   SIGNAL n2164 : STD_LOGIC;
   SIGNAL n2165 : STD_LOGIC;
   SIGNAL n2166 : STD_LOGIC;
   SIGNAL n2167 : STD_LOGIC;
   SIGNAL n2168 : STD_LOGIC;
   SIGNAL n2169 : STD_LOGIC;
   SIGNAL n2170 : STD_LOGIC;
   SIGNAL n2171 : STD_LOGIC;
   SIGNAL n2172 : STD_LOGIC;
   SIGNAL n2173 : STD_LOGIC;
   SIGNAL n2174 : STD_LOGIC;
   SIGNAL n2175 : STD_LOGIC;
   SIGNAL n2176 : STD_LOGIC;
   SIGNAL n2177 : STD_LOGIC;
   SIGNAL n2178 : STD_LOGIC;
   SIGNAL n2179 : STD_LOGIC;
   SIGNAL n2180 : STD_LOGIC;
   SIGNAL n2181 : STD_LOGIC;
   SIGNAL n2182 : STD_LOGIC;
   SIGNAL n2184 : STD_LOGIC;
   SIGNAL n2187 : STD_LOGIC;
   SIGNAL n2193 : STD_LOGIC;
   SIGNAL n2195 : STD_LOGIC;
   SIGNAL n2602 : STD_LOGIC;
   SIGNAL n2603 : STD_LOGIC;
   SIGNAL n2604 : STD_LOGIC;
   SIGNAL n2605 : STD_LOGIC;
   SIGNAL n2606 : STD_LOGIC;
   SIGNAL n2607 : STD_LOGIC;
   SIGNAL n2608 : STD_LOGIC;
   SIGNAL n2609 : STD_LOGIC;
   SIGNAL n2610 : STD_LOGIC;
   SIGNAL n2611 : STD_LOGIC;
   SIGNAL n2612 : STD_LOGIC;
   SIGNAL n2613 : STD_LOGIC;
   SIGNAL n2614 : STD_LOGIC;
   SIGNAL n2615 : STD_LOGIC;
   SIGNAL n2616 : STD_LOGIC;
   SIGNAL n2617 : STD_LOGIC;
   SIGNAL n2618 : STD_LOGIC;
   SIGNAL n2619 : STD_LOGIC;
   SIGNAL n2620 : STD_LOGIC;
   SIGNAL n2621 : STD_LOGIC;
   SIGNAL n2622 : STD_LOGIC;
   SIGNAL n2623 : STD_LOGIC;
   SIGNAL n2624 : STD_LOGIC;
   SIGNAL n2625 : STD_LOGIC;
   SIGNAL n2626 : STD_LOGIC;
   SIGNAL n2627 : STD_LOGIC;
   SIGNAL n2628 : STD_LOGIC;
   SIGNAL n2629 : STD_LOGIC;
   SIGNAL n2630 : STD_LOGIC;
   SIGNAL n2631 : STD_LOGIC;
   SIGNAL n2632 : STD_LOGIC;
   SIGNAL n2633 : STD_LOGIC;
   SIGNAL n2634 : STD_LOGIC;
   SIGNAL n2635 : STD_LOGIC;
   SIGNAL n2636 : STD_LOGIC;
   SIGNAL n2637 : STD_LOGIC;
   SIGNAL n2638 : STD_LOGIC;
   SIGNAL n2639 : STD_LOGIC;
   SIGNAL n2640 : STD_LOGIC;
   SIGNAL n2641 : STD_LOGIC;
   SIGNAL n2642 : STD_LOGIC;
   SIGNAL n2643 : STD_LOGIC;
   SIGNAL n2644 : STD_LOGIC;
   SIGNAL n2645 : STD_LOGIC;
   SIGNAL n2646 : STD_LOGIC;
   SIGNAL n2647 : STD_LOGIC;
   SIGNAL n2648 : STD_LOGIC;
   SIGNAL n2649 : STD_LOGIC;
   SIGNAL n2650 : STD_LOGIC;
   SIGNAL n2651 : STD_LOGIC;
   SIGNAL n2652 : STD_LOGIC;
   SIGNAL n2653 : STD_LOGIC;
   SIGNAL n2654 : STD_LOGIC;
   SIGNAL n2655 : STD_LOGIC;
   SIGNAL n2656 : STD_LOGIC;
   SIGNAL n2657 : STD_LOGIC;
   SIGNAL n2658 : STD_LOGIC;
   SIGNAL n2659 : STD_LOGIC;
   SIGNAL n2660 : STD_LOGIC;
   SIGNAL n2661 : STD_LOGIC;
   SIGNAL n2662 : STD_LOGIC;
   SIGNAL n2663 : STD_LOGIC;
   SIGNAL n2664 : STD_LOGIC;
   SIGNAL n2665 : STD_LOGIC;
   SIGNAL n2666 : STD_LOGIC;
   SIGNAL n2667 : STD_LOGIC;
   SIGNAL n2668 : STD_LOGIC;
   SIGNAL n2669 : STD_LOGIC;
   SIGNAL n2670 : STD_LOGIC;
   SIGNAL n2671 : STD_LOGIC;
   SIGNAL n2672 : STD_LOGIC;
   SIGNAL n2673 : STD_LOGIC;
   SIGNAL n2674 : STD_LOGIC;
   SIGNAL n2675 : STD_LOGIC;
   SIGNAL n2676 : STD_LOGIC;
   SIGNAL n2677 : STD_LOGIC;
   SIGNAL n2678 : STD_LOGIC;
   SIGNAL n2679 : STD_LOGIC;
   SIGNAL n2680 : STD_LOGIC;
   SIGNAL n2681 : STD_LOGIC;
   SIGNAL n2682 : STD_LOGIC;
   SIGNAL n2683 : STD_LOGIC;
   SIGNAL n2684 : STD_LOGIC;
   SIGNAL n2685 : STD_LOGIC;
   SIGNAL n2686 : STD_LOGIC;
   SIGNAL n2687 : STD_LOGIC;
   SIGNAL n2688 : STD_LOGIC;
   SIGNAL n2689 : STD_LOGIC;
   SIGNAL n2690 : STD_LOGIC;
   SIGNAL n2691 : STD_LOGIC;
   SIGNAL n2692 : STD_LOGIC;
   SIGNAL n2693 : STD_LOGIC;
   SIGNAL n2694 : STD_LOGIC;
   SIGNAL n2695 : STD_LOGIC;
   SIGNAL n2696 : STD_LOGIC;
   SIGNAL n2697 : STD_LOGIC;
   SIGNAL n2698 : STD_LOGIC;
   SIGNAL n2699 : STD_LOGIC;
   SIGNAL n2700 : STD_LOGIC;
   SIGNAL n2701 : STD_LOGIC;
   SIGNAL n2702 : STD_LOGIC;
   SIGNAL n2703 : STD_LOGIC;
   SIGNAL n2704 : STD_LOGIC;
   SIGNAL n2705 : STD_LOGIC;
   SIGNAL n2706 : STD_LOGIC;
   SIGNAL n2707 : STD_LOGIC;
   SIGNAL n2708 : STD_LOGIC;
   SIGNAL n2709 : STD_LOGIC;
   SIGNAL n2710 : STD_LOGIC;
   SIGNAL n2711 : STD_LOGIC;
   SIGNAL n2712 : STD_LOGIC;
   SIGNAL n2713 : STD_LOGIC;
   SIGNAL n2714 : STD_LOGIC;
   SIGNAL n2715 : STD_LOGIC;
   SIGNAL n2716 : STD_LOGIC;
   SIGNAL n2717 : STD_LOGIC;
   SIGNAL n2718 : STD_LOGIC;
   SIGNAL n2719 : STD_LOGIC;
   SIGNAL n2720 : STD_LOGIC;
   SIGNAL n2721 : STD_LOGIC;
   SIGNAL n2722 : STD_LOGIC;
   SIGNAL n2723 : STD_LOGIC;
   SIGNAL n2724 : STD_LOGIC;
   SIGNAL n2725 : STD_LOGIC;
   SIGNAL n2726 : STD_LOGIC;
   SIGNAL n2727 : STD_LOGIC;
   SIGNAL n2728 : STD_LOGIC;
   SIGNAL n2729 : STD_LOGIC;
   SIGNAL n2730 : STD_LOGIC;
   SIGNAL n2731 : STD_LOGIC;
   SIGNAL n2732 : STD_LOGIC;
   SIGNAL n2733 : STD_LOGIC;
   SIGNAL n2734 : STD_LOGIC;
   SIGNAL n2735 : STD_LOGIC;
   SIGNAL n2736 : STD_LOGIC;
   SIGNAL n2737 : STD_LOGIC;
   SIGNAL n2738 : STD_LOGIC;
   SIGNAL n2739 : STD_LOGIC;
   SIGNAL n2740 : STD_LOGIC;
   SIGNAL n2741 : STD_LOGIC;
   SIGNAL n2742 : STD_LOGIC;
   SIGNAL n2743 : STD_LOGIC;
   SIGNAL n2744 : STD_LOGIC;
   SIGNAL n2745 : STD_LOGIC;
   SIGNAL n2746 : STD_LOGIC;
   SIGNAL n2747 : STD_LOGIC;
   SIGNAL n2748 : STD_LOGIC;
   SIGNAL n2749 : STD_LOGIC;
   SIGNAL n2750 : STD_LOGIC;
   SIGNAL n2751 : STD_LOGIC;
   SIGNAL n2752 : STD_LOGIC;
   SIGNAL n2753 : STD_LOGIC;
   SIGNAL n2754 : STD_LOGIC;
   SIGNAL n2755 : STD_LOGIC;
   SIGNAL n2756 : STD_LOGIC;
   SIGNAL n2915 : STD_LOGIC;
   SIGNAL n2916 : STD_LOGIC;
   SIGNAL n2917 : STD_LOGIC;
   SIGNAL n2918 : STD_LOGIC;
   SIGNAL n2919 : STD_LOGIC;
   SIGNAL n2920 : STD_LOGIC;
   SIGNAL n2921 : STD_LOGIC;
   SIGNAL n2922 : STD_LOGIC;
   SIGNAL n2923 : STD_LOGIC;
   SIGNAL n2924 : STD_LOGIC;
   SIGNAL n2925 : STD_LOGIC;
   SIGNAL n2926 : STD_LOGIC;
   SIGNAL n2927 : STD_LOGIC;
   SIGNAL n2928 : STD_LOGIC;
   SIGNAL n2929 : STD_LOGIC;
   SIGNAL n2930 : STD_LOGIC;
   SIGNAL n2931 : STD_LOGIC;
   SIGNAL n2932 : STD_LOGIC;
   SIGNAL n2933 : STD_LOGIC;
   SIGNAL n2934 : STD_LOGIC;
   SIGNAL n2935 : STD_LOGIC;
   SIGNAL n2936 : STD_LOGIC;
   SIGNAL n2937 : STD_LOGIC;
   SIGNAL n2938 : STD_LOGIC;
   SIGNAL n2940 : STD_LOGIC;
   SIGNAL n2943 : STD_LOGIC;
   SIGNAL n2960 : STD_LOGIC;
   SIGNAL n2962 : STD_LOGIC;
   SIGNAL n3403 : STD_LOGIC;
   SIGNAL n3404 : STD_LOGIC;
   SIGNAL n3405 : STD_LOGIC;
   SIGNAL n3406 : STD_LOGIC;
   SIGNAL n3407 : STD_LOGIC;
   SIGNAL n3408 : STD_LOGIC;
   SIGNAL n3409 : STD_LOGIC;
   SIGNAL n3410 : STD_LOGIC;
   SIGNAL n3411 : STD_LOGIC;
   SIGNAL n3412 : STD_LOGIC;
   SIGNAL n3413 : STD_LOGIC;
   SIGNAL n3414 : STD_LOGIC;
   SIGNAL n3415 : STD_LOGIC;
   SIGNAL n3416 : STD_LOGIC;
   SIGNAL n3417 : STD_LOGIC;
   SIGNAL n3418 : STD_LOGIC;
   SIGNAL n3419 : STD_LOGIC;
   SIGNAL n3420 : STD_LOGIC;
   SIGNAL n3421 : STD_LOGIC;
   SIGNAL n3422 : STD_LOGIC;
   SIGNAL n3423 : STD_LOGIC;
   SIGNAL n3424 : STD_LOGIC;
   SIGNAL n3425 : STD_LOGIC;
   SIGNAL n3426 : STD_LOGIC;
   SIGNAL n3428 : STD_LOGIC;
   SIGNAL n3431 : STD_LOGIC;
   SIGNAL n3448 : STD_LOGIC;
   SIGNAL n3450 : STD_LOGIC;
   SIGNAL n4288 : STD_LOGIC;
   SIGNAL n6210 : STD_LOGIC;
   SIGNAL n6211 : STD_LOGIC;
   SIGNAL n6212 : STD_LOGIC;
   SIGNAL n6213 : STD_LOGIC;
   SIGNAL n6214 : STD_LOGIC;
   SIGNAL n6215 : STD_LOGIC;
   SIGNAL n6216 : STD_LOGIC;
   SIGNAL n6217 : STD_LOGIC;
   SIGNAL n6218 : STD_LOGIC;
   SIGNAL n6219 : STD_LOGIC;
   SIGNAL n6220 : STD_LOGIC;
   SIGNAL n6221 : STD_LOGIC;
   SIGNAL n6222 : STD_LOGIC;
   SIGNAL n6223 : STD_LOGIC;
   SIGNAL n6224 : STD_LOGIC;
   SIGNAL n6225 : STD_LOGIC;
   SIGNAL n6226 : STD_LOGIC;
   SIGNAL n6227 : STD_LOGIC;
   SIGNAL n6228 : STD_LOGIC;
   SIGNAL n6229 : STD_LOGIC;
   SIGNAL n6230 : STD_LOGIC;
   SIGNAL n6231 : STD_LOGIC;
   SIGNAL n6232 : STD_LOGIC;
   SIGNAL n6233 : STD_LOGIC;
   SIGNAL n6234 : STD_LOGIC;
   SIGNAL n6235 : STD_LOGIC;
   SIGNAL n6236 : STD_LOGIC;
   SIGNAL n6237 : STD_LOGIC;
   SIGNAL n6238 : STD_LOGIC;
   SIGNAL n6239 : STD_LOGIC;
   SIGNAL n6240 : STD_LOGIC;
   SIGNAL n6241 : STD_LOGIC;
   SIGNAL n6242 : STD_LOGIC;
   SIGNAL n6243 : STD_LOGIC;
   SIGNAL n6244 : STD_LOGIC;
   SIGNAL n6245 : STD_LOGIC;
   SIGNAL n6246 : STD_LOGIC;
   SIGNAL n6247 : STD_LOGIC;
   SIGNAL n6248 : STD_LOGIC;
   SIGNAL n6249 : STD_LOGIC;
   SIGNAL n6250 : STD_LOGIC;
   SIGNAL n6251 : STD_LOGIC;
   SIGNAL n6252 : STD_LOGIC;
   SIGNAL n6385 : STD_LOGIC;
   SIGNAL n6386 : STD_LOGIC;
   SIGNAL n6387 : STD_LOGIC;
   SIGNAL n6388 : STD_LOGIC;
   SIGNAL n6389 : STD_LOGIC;
   SIGNAL n6390 : STD_LOGIC;
   SIGNAL n6391 : STD_LOGIC;
   SIGNAL n6392 : STD_LOGIC;
   SIGNAL n6393 : STD_LOGIC;
   SIGNAL n6394 : STD_LOGIC;
   SIGNAL n6395 : STD_LOGIC;
   SIGNAL n6396 : STD_LOGIC;
   SIGNAL n6397 : STD_LOGIC;
   SIGNAL n6398 : STD_LOGIC;
   SIGNAL n6399 : STD_LOGIC;
   SIGNAL n6400 : STD_LOGIC;
   SIGNAL n6402 : STD_LOGIC;
   SIGNAL n6405 : STD_LOGIC;
   SIGNAL n6432 : STD_LOGIC;
   SIGNAL n6434 : STD_LOGIC;
   SIGNAL n6936 : STD_LOGIC;
   SIGNAL n6937 : STD_LOGIC;
   SIGNAL n6938 : STD_LOGIC;
   SIGNAL n6939 : STD_LOGIC;
   SIGNAL n6940 : STD_LOGIC;
   SIGNAL n6941 : STD_LOGIC;
   SIGNAL n6942 : STD_LOGIC;
   SIGNAL n6943 : STD_LOGIC;
   SIGNAL n6944 : STD_LOGIC;
   SIGNAL n6945 : STD_LOGIC;
   SIGNAL n6946 : STD_LOGIC;
   SIGNAL n6947 : STD_LOGIC;
   SIGNAL n6948 : STD_LOGIC;
   SIGNAL n6949 : STD_LOGIC;
   SIGNAL n6950 : STD_LOGIC;
   SIGNAL n6951 : STD_LOGIC;
   SIGNAL n6952 : STD_LOGIC;
   SIGNAL n6953 : STD_LOGIC;
   SIGNAL n6954 : STD_LOGIC;
   SIGNAL n6955 : STD_LOGIC;
   SIGNAL n6956 : STD_LOGIC;
   SIGNAL n6957 : STD_LOGIC;
   SIGNAL n6958 : STD_LOGIC;
   SIGNAL n6959 : STD_LOGIC;
   SIGNAL n6960 : STD_LOGIC;
   SIGNAL n6961 : STD_LOGIC;
   SIGNAL n6962 : STD_LOGIC;
   SIGNAL n6963 : STD_LOGIC;
   SIGNAL n6964 : STD_LOGIC;
   SIGNAL n6965 : STD_LOGIC;
   SIGNAL n6967 : STD_LOGIC;
   SIGNAL n6970 : STD_LOGIC;
   SIGNAL n6975 : STD_LOGIC;
   SIGNAL n6977 : STD_LOGIC;
   SIGNAL n7477 : STD_LOGIC;
   SIGNAL n7478 : STD_LOGIC;
   SIGNAL n7479 : STD_LOGIC;
   SIGNAL n7480 : STD_LOGIC;
   SIGNAL n7481 : STD_LOGIC;
   SIGNAL n7482 : STD_LOGIC;
   SIGNAL n7483 : STD_LOGIC;
   SIGNAL n7484 : STD_LOGIC;
   SIGNAL n7485 : STD_LOGIC;
   SIGNAL n7486 : STD_LOGIC;
   SIGNAL n7487 : STD_LOGIC;
   SIGNAL n7488 : STD_LOGIC;
   SIGNAL n7489 : STD_LOGIC;
   SIGNAL n7490 : STD_LOGIC;
   SIGNAL n7491 : STD_LOGIC;
   SIGNAL n7492 : STD_LOGIC;
   SIGNAL n7493 : STD_LOGIC;
   SIGNAL n7494 : STD_LOGIC;
   SIGNAL n7495 : STD_LOGIC;
   SIGNAL n7496 : STD_LOGIC;
   SIGNAL n7497 : STD_LOGIC;
   SIGNAL n7498 : STD_LOGIC;
   SIGNAL n7499 : STD_LOGIC;
   SIGNAL n7500 : STD_LOGIC;
   SIGNAL n7501 : STD_LOGIC;
   SIGNAL n7502 : STD_LOGIC;
   SIGNAL n7503 : STD_LOGIC;
   SIGNAL n7504 : STD_LOGIC;
   SIGNAL n7505 : STD_LOGIC;
   SIGNAL n7506 : STD_LOGIC;
   SIGNAL n7508 : STD_LOGIC;
   SIGNAL n7511 : STD_LOGIC;
   SIGNAL n7516 : STD_LOGIC;
   SIGNAL n7518 : STD_LOGIC;

BEGIN

   n135 <= DIN(0);
   n136 <= DIN(1);
   n137 <= DIN(2);
   n138 <= DIN(3);
   n139 <= DIN(4);
   n140 <= DIN(5);
   n141 <= DIN(6);
   n142 <= DIN(7);
   n143 <= DIN(8);
   n144 <= DIN(9);
   n145 <= DIN(10);
   n146 <= DIN(11);
   n147 <= DIN(12);
   n148 <= DIN(13);
   n149 <= ND;
   n152 <= CLK;
   n153 <= ADDR(0);
   n154 <= ADDR(1);
   n155 <= ADDR(2);
   n156 <= ADDR(3);
   n157 <= ADDR(4);
   n158 <= LD_DIN(0);
   n159 <= LD_DIN(1);
   n160 <= LD_DIN(2);
   n161 <= LD_DIN(3);
   n162 <= LD_DIN(4);
   n163 <= LD_DIN(5);
   n164 <= LD_DIN(6);
   n165 <= LD_DIN(7);
   n166 <= LD_DIN(8);
   n167 <= LD_DIN(9);
   n168 <= LD_DIN(10);
   n169 <= LD_DIN(11);
   n170 <= LD_DIN(12);
   n171 <= LD_DIN(13);
   n172 <= LD_DIN(14);
   n173 <= LD_DIN(15);
   n174 <= LD_DIN(16);
   n175 <= LD_DIN(17);
   n176 <= LD_DIN(18);
   n177 <= LD_DIN(19);
   n178 <= LD_DIN(20);
   n179 <= LD_DIN(21);
   n180 <= LD_DIN(22);
   n181 <= LD_DIN(23);
   n182 <= LD_DIN(24);
   n183 <= LD_DIN(25);
   n184 <= LD_DIN(26);
   n185 <= LD_DIN(27);
   n186 <= LD_DIN(28);
   n187 <= LD_DIN(29);
   n188 <= LD_DIN(30);
   n189 <= LD_DIN(31);
   n190 <= WE;
   n191 <= SEL;
   RDY <= n150;
   RFD <= n151;
   DOUT_I(0) <= n192;
   DOUT_I(1) <= n193;
   DOUT_I(2) <= n194;
   DOUT_I(3) <= n195;
   DOUT_I(4) <= n196;
   DOUT_I(5) <= n197;
   DOUT_I(6) <= n198;
   DOUT_I(7) <= n199;
   DOUT_I(8) <= n200;
   DOUT_I(9) <= n201;
   DOUT_I(10) <= n202;
   DOUT_I(11) <= n203;
   DOUT_I(12) <= n204;
   DOUT_I(13) <= n205;
   DOUT_I(14) <= n206;
   DOUT_I(15) <= n207;
   DOUT_I(16) <= n208;
   DOUT_I(17) <= n209;
   DOUT_I(18) <= n210;
   DOUT_I(19) <= n211;
   DOUT_I(20) <= n212;
   DOUT_I(21) <= n213;
   DOUT_I(22) <= n214;
   DOUT_I(23) <= n215;
   DOUT_I(24) <= n216;
   DOUT_I(25) <= n217;
   DOUT_I(26) <= n218;
   DOUT_I(27) <= n219;
   DOUT_I(28) <= n220;
   DOUT_I(29) <= n221;
   DOUT_Q(0) <= n222;
   DOUT_Q(1) <= n223;
   DOUT_Q(2) <= n224;
   DOUT_Q(3) <= n225;
   DOUT_Q(4) <= n226;
   DOUT_Q(5) <= n227;
   DOUT_Q(6) <= n228;
   DOUT_Q(7) <= n229;
   DOUT_Q(8) <= n230;
   DOUT_Q(9) <= n231;
   DOUT_Q(10) <= n232;
   DOUT_Q(11) <= n233;
   DOUT_Q(12) <= n234;
   DOUT_Q(13) <= n235;
   DOUT_Q(14) <= n236;
   DOUT_Q(15) <= n237;
   DOUT_Q(16) <= n238;
   DOUT_Q(17) <= n239;
   DOUT_Q(18) <= n240;
   DOUT_Q(19) <= n241;
   DOUT_Q(20) <= n242;
   DOUT_Q(21) <= n243;
   DOUT_Q(22) <= n244;
   DOUT_Q(23) <= n245;
   DOUT_Q(24) <= n246;
   DOUT_Q(25) <= n247;
   DOUT_Q(26) <= n248;
   DOUT_Q(27) <= n249;
   DOUT_Q(28) <= n250;
   DOUT_Q(29) <= n251;

   BU4_I0 <= n157;
   BU4_I1 <= n156;
   BU4_I2 <= n155;
   BU4_I3 <= n191;
   n54 <= BU4_O;
   BU4 : LUT4
      GENERIC MAP (
         INIT  => X"1000"
      )
      PORT MAP (
         I0 => BU4_I0,
         I1 => BU4_I1,
         I2 => BU4_I2,
         I3 => BU4_I3,
         O => BU4_O
      );

   BU8_I0 <= n54;
   BU8_I1 <= n190;
   BU8_I2 <= n154;
   BU8_I3 <= n153;
   n291 <= BU8_O;
   BU8 : LUT4
      GENERIC MAP (
         INIT  => X"0080"
      )
      PORT MAP (
         I0 => BU8_I0,
         I1 => BU8_I1,
         I2 => BU8_I2,
         I3 => BU8_I3,
         O => BU8_O
      );

   BU10_I0 <= '1';
   BU10_I1 <= '0';
   BU10_I2 <= '0';
   BU10_I3 <= '0';
   n151 <= BU10_O;
   BU10 : LUT4
      GENERIC MAP (
         INIT  => X"aaaa"
      )
      PORT MAP (
         I0 => BU10_I0,
         I1 => BU10_I1,
         I2 => BU10_I2,
         I3 => BU10_I3,
         O => BU10_O
      );

   BU1292_D <= n149;
   BU1292_C <= n152;
   BU1292_CE <= '1';
   n340 <= BU1292_Q;
   BU1292 : FDE
      PORT MAP (
         D => BU1292_D,
         C => BU1292_C,
         CE => BU1292_CE,
         Q => BU1292_Q
      );

   BU14_D <= n135;
   BU14_CE <= n149;
   BU14_CLK <= n152;
   BU14_A0 <= '0';
   BU14_A1 <= '1';
   BU14_A2 <= '0';
   BU14_A3 <= '0';
   n924 <= BU14_Q;
   BU14 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU14_D,
         CE => BU14_CE,
         CLK => BU14_CLK,
         A0 => BU14_A0,
         A1 => BU14_A1,
         A2 => BU14_A2,
         A3 => BU14_A3,
         Q => BU14_Q
      );

   BU16_D <= n924;
   BU16_C <= n152;
   BU16_CE <= n149;
   n587 <= BU16_Q;
   BU16 : FDE
      PORT MAP (
         D => BU16_D,
         C => BU16_C,
         CE => BU16_CE,
         Q => BU16_Q
      );

   BU17_D <= n136;
   BU17_CE <= n149;
   BU17_CLK <= n152;
   BU17_A0 <= '0';
   BU17_A1 <= '1';
   BU17_A2 <= '0';
   BU17_A3 <= '0';
   n925 <= BU17_Q;
   BU17 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU17_D,
         CE => BU17_CE,
         CLK => BU17_CLK,
         A0 => BU17_A0,
         A1 => BU17_A1,
         A2 => BU17_A2,
         A3 => BU17_A3,
         Q => BU17_Q
      );

   BU19_D <= n925;
   BU19_C <= n152;
   BU19_CE <= n149;
   n586 <= BU19_Q;
   BU19 : FDE
      PORT MAP (
         D => BU19_D,
         C => BU19_C,
         CE => BU19_CE,
         Q => BU19_Q
      );

   BU20_D <= n137;
   BU20_CE <= n149;
   BU20_CLK <= n152;
   BU20_A0 <= '0';
   BU20_A1 <= '1';
   BU20_A2 <= '0';
   BU20_A3 <= '0';
   n926 <= BU20_Q;
   BU20 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU20_D,
         CE => BU20_CE,
         CLK => BU20_CLK,
         A0 => BU20_A0,
         A1 => BU20_A1,
         A2 => BU20_A2,
         A3 => BU20_A3,
         Q => BU20_Q
      );

   BU22_D <= n926;
   BU22_C <= n152;
   BU22_CE <= n149;
   n585 <= BU22_Q;
   BU22 : FDE
      PORT MAP (
         D => BU22_D,
         C => BU22_C,
         CE => BU22_CE,
         Q => BU22_Q
      );

   BU23_D <= n138;
   BU23_CE <= n149;
   BU23_CLK <= n152;
   BU23_A0 <= '0';
   BU23_A1 <= '1';
   BU23_A2 <= '0';
   BU23_A3 <= '0';
   n927 <= BU23_Q;
   BU23 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU23_D,
         CE => BU23_CE,
         CLK => BU23_CLK,
         A0 => BU23_A0,
         A1 => BU23_A1,
         A2 => BU23_A2,
         A3 => BU23_A3,
         Q => BU23_Q
      );

   BU25_D <= n927;
   BU25_C <= n152;
   BU25_CE <= n149;
   n584 <= BU25_Q;
   BU25 : FDE
      PORT MAP (
         D => BU25_D,
         C => BU25_C,
         CE => BU25_CE,
         Q => BU25_Q
      );

   BU26_D <= n139;
   BU26_CE <= n149;
   BU26_CLK <= n152;
   BU26_A0 <= '0';
   BU26_A1 <= '1';
   BU26_A2 <= '0';
   BU26_A3 <= '0';
   n928 <= BU26_Q;
   BU26 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU26_D,
         CE => BU26_CE,
         CLK => BU26_CLK,
         A0 => BU26_A0,
         A1 => BU26_A1,
         A2 => BU26_A2,
         A3 => BU26_A3,
         Q => BU26_Q
      );

   BU28_D <= n928;
   BU28_C <= n152;
   BU28_CE <= n149;
   n583 <= BU28_Q;
   BU28 : FDE
      PORT MAP (
         D => BU28_D,
         C => BU28_C,
         CE => BU28_CE,
         Q => BU28_Q
      );

   BU29_D <= n140;
   BU29_CE <= n149;
   BU29_CLK <= n152;
   BU29_A0 <= '0';
   BU29_A1 <= '1';
   BU29_A2 <= '0';
   BU29_A3 <= '0';
   n929 <= BU29_Q;
   BU29 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU29_D,
         CE => BU29_CE,
         CLK => BU29_CLK,
         A0 => BU29_A0,
         A1 => BU29_A1,
         A2 => BU29_A2,
         A3 => BU29_A3,
         Q => BU29_Q
      );

   BU31_D <= n929;
   BU31_C <= n152;
   BU31_CE <= n149;
   n582 <= BU31_Q;
   BU31 : FDE
      PORT MAP (
         D => BU31_D,
         C => BU31_C,
         CE => BU31_CE,
         Q => BU31_Q
      );

   BU32_D <= n141;
   BU32_CE <= n149;
   BU32_CLK <= n152;
   BU32_A0 <= '0';
   BU32_A1 <= '1';
   BU32_A2 <= '0';
   BU32_A3 <= '0';
   n930 <= BU32_Q;
   BU32 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU32_D,
         CE => BU32_CE,
         CLK => BU32_CLK,
         A0 => BU32_A0,
         A1 => BU32_A1,
         A2 => BU32_A2,
         A3 => BU32_A3,
         Q => BU32_Q
      );

   BU34_D <= n930;
   BU34_C <= n152;
   BU34_CE <= n149;
   n581 <= BU34_Q;
   BU34 : FDE
      PORT MAP (
         D => BU34_D,
         C => BU34_C,
         CE => BU34_CE,
         Q => BU34_Q
      );

   BU35_D <= n142;
   BU35_CE <= n149;
   BU35_CLK <= n152;
   BU35_A0 <= '0';
   BU35_A1 <= '1';
   BU35_A2 <= '0';
   BU35_A3 <= '0';
   n931 <= BU35_Q;
   BU35 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU35_D,
         CE => BU35_CE,
         CLK => BU35_CLK,
         A0 => BU35_A0,
         A1 => BU35_A1,
         A2 => BU35_A2,
         A3 => BU35_A3,
         Q => BU35_Q
      );

   BU37_D <= n931;
   BU37_C <= n152;
   BU37_CE <= n149;
   n580 <= BU37_Q;
   BU37 : FDE
      PORT MAP (
         D => BU37_D,
         C => BU37_C,
         CE => BU37_CE,
         Q => BU37_Q
      );

   BU38_D <= n143;
   BU38_CE <= n149;
   BU38_CLK <= n152;
   BU38_A0 <= '0';
   BU38_A1 <= '1';
   BU38_A2 <= '0';
   BU38_A3 <= '0';
   n932 <= BU38_Q;
   BU38 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU38_D,
         CE => BU38_CE,
         CLK => BU38_CLK,
         A0 => BU38_A0,
         A1 => BU38_A1,
         A2 => BU38_A2,
         A3 => BU38_A3,
         Q => BU38_Q
      );

   BU40_D <= n932;
   BU40_C <= n152;
   BU40_CE <= n149;
   n579 <= BU40_Q;
   BU40 : FDE
      PORT MAP (
         D => BU40_D,
         C => BU40_C,
         CE => BU40_CE,
         Q => BU40_Q
      );

   BU41_D <= n144;
   BU41_CE <= n149;
   BU41_CLK <= n152;
   BU41_A0 <= '0';
   BU41_A1 <= '1';
   BU41_A2 <= '0';
   BU41_A3 <= '0';
   n933 <= BU41_Q;
   BU41 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU41_D,
         CE => BU41_CE,
         CLK => BU41_CLK,
         A0 => BU41_A0,
         A1 => BU41_A1,
         A2 => BU41_A2,
         A3 => BU41_A3,
         Q => BU41_Q
      );

   BU43_D <= n933;
   BU43_C <= n152;
   BU43_CE <= n149;
   n578 <= BU43_Q;
   BU43 : FDE
      PORT MAP (
         D => BU43_D,
         C => BU43_C,
         CE => BU43_CE,
         Q => BU43_Q
      );

   BU44_D <= n145;
   BU44_CE <= n149;
   BU44_CLK <= n152;
   BU44_A0 <= '0';
   BU44_A1 <= '1';
   BU44_A2 <= '0';
   BU44_A3 <= '0';
   n934 <= BU44_Q;
   BU44 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU44_D,
         CE => BU44_CE,
         CLK => BU44_CLK,
         A0 => BU44_A0,
         A1 => BU44_A1,
         A2 => BU44_A2,
         A3 => BU44_A3,
         Q => BU44_Q
      );

   BU46_D <= n934;
   BU46_C <= n152;
   BU46_CE <= n149;
   n577 <= BU46_Q;
   BU46 : FDE
      PORT MAP (
         D => BU46_D,
         C => BU46_C,
         CE => BU46_CE,
         Q => BU46_Q
      );

   BU47_D <= n146;
   BU47_CE <= n149;
   BU47_CLK <= n152;
   BU47_A0 <= '0';
   BU47_A1 <= '1';
   BU47_A2 <= '0';
   BU47_A3 <= '0';
   n935 <= BU47_Q;
   BU47 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU47_D,
         CE => BU47_CE,
         CLK => BU47_CLK,
         A0 => BU47_A0,
         A1 => BU47_A1,
         A2 => BU47_A2,
         A3 => BU47_A3,
         Q => BU47_Q
      );

   BU49_D <= n935;
   BU49_C <= n152;
   BU49_CE <= n149;
   n576 <= BU49_Q;
   BU49 : FDE
      PORT MAP (
         D => BU49_D,
         C => BU49_C,
         CE => BU49_CE,
         Q => BU49_Q
      );

   BU50_D <= n147;
   BU50_CE <= n149;
   BU50_CLK <= n152;
   BU50_A0 <= '0';
   BU50_A1 <= '1';
   BU50_A2 <= '0';
   BU50_A3 <= '0';
   n936 <= BU50_Q;
   BU50 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU50_D,
         CE => BU50_CE,
         CLK => BU50_CLK,
         A0 => BU50_A0,
         A1 => BU50_A1,
         A2 => BU50_A2,
         A3 => BU50_A3,
         Q => BU50_Q
      );

   BU52_D <= n936;
   BU52_C <= n152;
   BU52_CE <= n149;
   n575 <= BU52_Q;
   BU52 : FDE
      PORT MAP (
         D => BU52_D,
         C => BU52_C,
         CE => BU52_CE,
         Q => BU52_Q
      );

   BU53_D <= n148;
   BU53_CE <= n149;
   BU53_CLK <= n152;
   BU53_A0 <= '0';
   BU53_A1 <= '1';
   BU53_A2 <= '0';
   BU53_A3 <= '0';
   n937 <= BU53_Q;
   BU53 : SRL16E
      GENERIC MAP (
         INIT  => X"0000"
      )
      PORT MAP (
         D => BU53_D,
         CE => BU53_CE,
         CLK => BU53_CLK,
         A0 => BU53_A0,
         A1 => BU53_A1,
         A2 => BU53_A2,
         A3 => BU53_A3,
         Q => BU53_Q
      );

   BU55_D <= n937;
   BU55_C <= n152;
   BU55_CE <= n149;
   n574 <= BU55_Q;
   BU55 : FDE
      PORT MAP (
         D => BU55_D,
         C => BU55_C,
         CE => BU55_CE,
         Q => BU55_Q
      );

   BU57_DATA(0) <= n158;
   BU57_DATA(1) <= n159;
   BU57_DATA(2) <= n160;
   BU57_DATA(3) <= n161;
   BU57_DATA(4) <= n162;
   BU57_DATA(5) <= n163;
   BU57_DATA(6) <= n164;
   BU57_DATA(7) <= n165;
   BU57_DATA(8) <= n166;
   BU57_DATA(9) <= n167;
   BU57_DATA(10) <= n168;
   BU57_DATA(11) <= n169;
   BU57_DATA(12) <= n170;
   BU57_DATA(13) <= n171;
   BU57_DATA(14) <= n172;
   BU57_DATA(15) <= n173;
   BU57_DATA(16) <= n174;
   BU57_DATA(17) <= n175;
   BU57_DATA(18) <= n176;
   BU57_DATA(19) <= n177;
   BU57_DATA(20) <= n178;
   BU57_DATA(21) <= n179;
   BU57_DATA(22) <= n180;
   BU57_DATA(23) <= n181;
   BU57_DATA(24) <= n182;
   BU57_DATA(25) <= n183;
   BU57_DATA(26) <= n184;
   BU57_DATA(27) <= n185;
   BU57_DATA(28) <= n186;
   BU57_DATA(29) <= n187;
   BU57_DATA(30) <= n188;
   BU57_DATA(31) <= n189;
   BU57_WE <= n291;
   BU57_CLK <= n152;
   BU57_CE <= n149;
   n339 <= BU57_RDY;
   n426 <= BU57_SINE(0);
   n425 <= BU57_SINE(1);
   n424 <= BU57_SINE(2);
   n423 <= BU57_SINE(3);
   n422 <= BU57_SINE(4);
   n421 <= BU57_SINE(5);
   n420 <= BU57_SINE(6);
   n419 <= BU57_SINE(7);
   n418 <= BU57_SINE(8);
   n417 <= BU57_SINE(9);
   n416 <= BU57_SINE(10);
   n415 <= BU57_SINE(11);
   n414 <= BU57_SINE(12);
   n413 <= BU57_SINE(13);
   n412 <= BU57_SINE(14);
   n630 <= BU57_COSINE(0);
   n629 <= BU57_COSINE(1);
   n628 <= BU57_COSINE(2);
   n627 <= BU57_COSINE(3);
   n626 <= BU57_COSINE(4);
   n625 <= BU57_COSINE(5);
   n624 <= BU57_COSINE(6);
   n623 <= BU57_COSINE(7);
   n622 <= BU57_COSINE(8);
   n621 <= BU57_COSINE(9);
   n620 <= BU57_COSINE(10);
   n619 <= BU57_COSINE(11);
   n618 <= BU57_COSINE(12);
   n617 <= BU57_COSINE(13);
   n616 <= BU57_COSINE(14);
   BU57 : C_DDS_V4_1
      GENERIC MAP (
         c_phase_offset_value => "00000000000000000000000000000000",
         c_phase_increment_value => "01001100110011001100110011001101",
         c_has_rdy => 1,
         c_has_sclr => 0,
         c_phase_offset => 0,
         c_data_width => 32,
         c_accumulator_latency => 1,
         c_enable_rlocs => 0,
         c_phase_angle_width => 13,
         c_has_rfd => 0,
         c_phase_increment => 1,
         c_negative_sine => 0,
         c_latency => 4,
         c_has_ce => 1,
         c_has_aclr => 0,
         c_outputs_required => 2,
         c_pipelined => 1,
         c_accumulator_width => 32,
         c_mem_type => 1,
         c_negative_cosine => 0,
         c_noise_shaping => 1,
         c_output_width => 15
      )
      PORT MAP (
         DATA => BU57_DATA,
         WE => BU57_WE,
         CLK => BU57_CLK,
         CE => BU57_CE,
         RDY => BU57_RDY,
         SINE => BU57_SINE,
         COSINE => BU57_COSINE
      );

   BU1294_I0 <= n339;
   BU1294_I1 <= n340;
   BU1294_I2 <= '0';
   BU1294_I3 <= '0';
   n338 <= BU1294_O;
   BU1294 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU1294_I0,
         I1 => BU1294_I1,
         I2 => BU1294_I2,
         I3 => BU1294_I3,
         O => BU1294_O
      );

   BU1296_clk <= n152;
   BU1296_a(13) <= n574;
   BU1296_a(12) <= n575;
   BU1296_a(11) <= n576;
   BU1296_a(10) <= n577;
   BU1296_a(9) <= n578;
   BU1296_a(8) <= n579;
   BU1296_a(7) <= n580;
   BU1296_a(6) <= n581;
   BU1296_a(5) <= n582;
   BU1296_a(4) <= n583;
   BU1296_a(3) <= n584;
   BU1296_a(2) <= n585;
   BU1296_a(1) <= n586;
   BU1296_a(0) <= n587;
   BU1296_b(14) <= n412;
   BU1296_b(13) <= n413;
   BU1296_b(12) <= n414;
   BU1296_b(11) <= n415;
   BU1296_b(10) <= n416;
   BU1296_b(9) <= n417;
   BU1296_b(8) <= n418;
   BU1296_b(7) <= n419;
   BU1296_b(6) <= n420;
   BU1296_b(5) <= n421;
   BU1296_b(4) <= n422;
   BU1296_b(3) <= n423;
   BU1296_b(2) <= n424;
   BU1296_b(1) <= n425;
   BU1296_b(0) <= n426;
   n457 <= BU1296_q(28);
   n458 <= BU1296_q(27);
   n459 <= BU1296_q(26);
   n460 <= BU1296_q(25);
   n461 <= BU1296_q(24);
   n462 <= BU1296_q(23);
   n463 <= BU1296_q(22);
   n464 <= BU1296_q(21);
   n465 <= BU1296_q(20);
   n466 <= BU1296_q(19);
   n467 <= BU1296_q(18);
   n468 <= BU1296_q(17);
   n469 <= BU1296_q(16);
   n470 <= BU1296_q(15);
   n471 <= BU1296_q(14);
   n472 <= BU1296_q(13);
   n473 <= BU1296_q(12);
   n474 <= BU1296_q(11);
   n475 <= BU1296_q(10);
   n476 <= BU1296_q(9);
   n477 <= BU1296_q(8);
   n478 <= BU1296_q(7);
   n479 <= BU1296_q(6);
   n480 <= BU1296_q(5);
   n481 <= BU1296_q(4);
   n482 <= BU1296_q(3);
   n483 <= BU1296_q(2);
   n484 <= BU1296_q(1);
   n485 <= BU1296_q(0);
   BU1296_a_signed <= '0';
   BU1296_loadb <= '0';
   BU1296_swapb <= '0';
   BU1296_ce <= '1';
   BU1296_aclr <= '0';
   BU1296_sclr <= '0';
   BU1296_nd <= n338;
   n544 <= BU1296_rdy;
   BU1296 : mult_gen_v5_0
      GENERIC MAP (
         c_a_width => 14,
         c_out_width => 29,
         c_b_type => 0,
         c_has_b => 1,
         c_has_rdy => 1,
         bram_addr_width => 8,
         c_has_sclr => 0,
         c_has_nd => 1,
         c_reg_a_b_inputs => 1,
         c_enable_rlocs => 0,
         c_has_rfd => 1,
         c_mult_type => 1,
         c_has_swapb => 0,
         c_baat => 14,
         c_use_luts => 1,
         c_has_load_done => 0,
         c_has_a_signed => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 1,
         c_output_hold => 0,
         c_stack_adders => 0,
         c_mem_type => 0,
         c_b_constant => 0,
         c_has_q => 1,
         c_has_loadb => 0,
         c_pipeline => 1,
         c_has_o => 0,
         c_standalone => 1,
         c_mem_init_prefix => "mem",
         c_a_type => 0,
         c_b_width => 15,
         c_sqm_type => 0,
         c_b_value => "0"
      )
      PORT MAP (
         clk => BU1296_clk,
         a => BU1296_a,
         b => BU1296_b,
         o => BU1296_o,
         q => BU1296_q,
         a_signed => BU1296_a_signed,
         loadb => BU1296_loadb,
         load_done => BU1296_load_done,
         swapb => BU1296_swapb,
         ce => BU1296_ce,
         aclr => BU1296_aclr,
         sclr => BU1296_sclr,
         rfd => BU1296_rfd,
         nd => BU1296_nd,
         rdy => BU1296_rdy
      );

   BU1517_I(0) <= n485;
   BU1517_I(1) <= n484;
   BU1517_I(2) <= n483;
   BU1517_I(3) <= n482;
   BU1517_I(4) <= n481;
   n1544 <= BU1517_O;
   BU1517 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 5,
         c_input_inv_mask => "01111"
      )
      PORT MAP (
         I => BU1517_I,
         O => BU1517_O
      );

   BU1526_I0 <= n480;
   BU1526_I1 <= n481;
   BU1526_I2 <= n1544;
   BU1526_I3 <= '0';
   n1541 <= BU1526_O;
   BU1526 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU1526_I0,
         I1 => BU1526_I1,
         I2 => BU1526_I2,
         I3 => BU1526_I3,
         O => BU1526_O
      );

   BU1527_A(0) <= n480;
   BU1527_A(1) <= n479;
   BU1527_A(2) <= n478;
   BU1527_A(3) <= n477;
   BU1527_A(4) <= n476;
   BU1527_A(5) <= n475;
   BU1527_A(6) <= n474;
   BU1527_A(7) <= n473;
   BU1527_A(8) <= n472;
   BU1527_A(9) <= n471;
   BU1527_A(10) <= n470;
   BU1527_A(11) <= n469;
   BU1527_A(12) <= n468;
   BU1527_A(13) <= n467;
   BU1527_A(14) <= n466;
   BU1527_A(15) <= n465;
   BU1527_A(16) <= n464;
   BU1527_A(17) <= n463;
   BU1527_A(18) <= n462;
   BU1527_A(19) <= n461;
   BU1527_A(20) <= n460;
   BU1527_A(21) <= n459;
   BU1527_A(22) <= n458;
   BU1527_A(23) <= n457;
   BU1527_B(0) <= n1541;
   n1516 <= BU1527_S(0);
   n1517 <= BU1527_S(1);
   n1518 <= BU1527_S(2);
   n1519 <= BU1527_S(3);
   n1520 <= BU1527_S(4);
   n1521 <= BU1527_S(5);
   n1522 <= BU1527_S(6);
   n1523 <= BU1527_S(7);
   n1524 <= BU1527_S(8);
   n1525 <= BU1527_S(9);
   n1526 <= BU1527_S(10);
   n1527 <= BU1527_S(11);
   n1528 <= BU1527_S(12);
   n1529 <= BU1527_S(13);
   n1530 <= BU1527_S(14);
   n1531 <= BU1527_S(15);
   n1532 <= BU1527_S(16);
   n1533 <= BU1527_S(17);
   n1534 <= BU1527_S(18);
   n1535 <= BU1527_S(19);
   n1536 <= BU1527_S(20);
   n1537 <= BU1527_S(21);
   n1538 <= BU1527_S(22);
   n1539 <= BU1527_S(23);
   BU1527 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU1527_A,
         B => BU1527_B,
         S => BU1527_S
      );

   BU1628_I0 <= n457;
   BU1628_I1 <= n458;
   BU1628_I2 <= n1539;
   BU1628_I3 <= '0';
   n1550 <= BU1628_O;
   BU1628 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU1628_I0,
         I1 => BU1628_I1,
         I2 => BU1628_I2,
         I3 => BU1628_I3,
         O => BU1628_O
      );

   BU1630_I0 <= n457;
   BU1630_I1 <= n1539;
   BU1630_I2 <= '0';
   BU1630_I3 <= '0';
   n1552 <= BU1630_O;
   BU1630 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU1630_I0,
         I1 => BU1630_I1,
         I2 => BU1630_I2,
         I3 => BU1630_I3,
         O => BU1630_O
      );

   BU1631_D(0) <= n1516;
   BU1631_D(1) <= n1517;
   BU1631_D(2) <= n1518;
   BU1631_D(3) <= n1519;
   BU1631_D(4) <= n1520;
   BU1631_D(5) <= n1521;
   BU1631_D(6) <= n1522;
   BU1631_D(7) <= n1523;
   BU1631_D(8) <= n1524;
   BU1631_D(9) <= n1525;
   BU1631_D(10) <= n1526;
   BU1631_D(11) <= n1527;
   BU1631_D(12) <= n1528;
   BU1631_D(13) <= n1529;
   BU1631_D(14) <= n1530;
   BU1631_D(15) <= n1531;
   BU1631_D(16) <= n1532;
   BU1631_D(17) <= n1533;
   BU1631_D(18) <= n1534;
   BU1631_D(19) <= n1535;
   BU1631_D(20) <= n1536;
   BU1631_D(21) <= n1537;
   BU1631_D(22) <= n1538;
   n3 <= BU1631_Q(0);
   n4 <= BU1631_Q(1);
   n5 <= BU1631_Q(2);
   n6 <= BU1631_Q(3);
   n7 <= BU1631_Q(4);
   n8 <= BU1631_Q(5);
   n9 <= BU1631_Q(6);
   n10 <= BU1631_Q(7);
   n11 <= BU1631_Q(8);
   n12 <= BU1631_Q(9);
   n13 <= BU1631_Q(10);
   n14 <= BU1631_Q(11);
   n15 <= BU1631_Q(12);
   n16 <= BU1631_Q(13);
   n17 <= BU1631_Q(14);
   n18 <= BU1631_Q(15);
   n19 <= BU1631_Q(16);
   n20 <= BU1631_Q(17);
   n21 <= BU1631_Q(18);
   n22 <= BU1631_Q(19);
   n23 <= BU1631_Q(20);
   n24 <= BU1631_Q(21);
   n25 <= BU1631_Q(22);
   BU1631_CLK <= n152;
   BU1631_SCLR <= n1550;
   BU1631_SSET <= n1552;
   BU1631 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU1631_D,
         Q => BU1631_Q,
         CLK => BU1631_CLK,
         SCLR => BU1631_SCLR,
         SSET => BU1631_SSET
      );

   BU1724_D(0) <= n1539;
   n26 <= BU1724_Q(0);
   BU1724_CLK <= n152;
   BU1724_SCLR <= n1552;
   BU1724_SSET <= n1550;
   BU1724 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU1724_D,
         Q => BU1724_Q,
         CLK => BU1724_CLK,
         SCLR => BU1724_SCLR,
         SSET => BU1724_SSET
      );

   BU1729_CLK <= n152;
   BU1729_D(0) <= n544;
   n2 <= BU1729_Q(0);
   BU1729 : C_SHIFT_RAM_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_read_mif => 0,
         c_has_a => 0,
         c_sync_priority => 0,
         c_has_sclr => 0,
         c_width => 1,
         c_enable_rlocs => 0,
         c_default_data_radix => 2,
         c_generate_mif => 0,
         c_ainit_val => "0",
         c_has_ce => 0,
         c_has_aclr => 0,
         c_mem_init_radix => 2,
         c_sync_enable => 0,
         c_depth => 1,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_shift_type => 0,
         c_mem_init_file => "null",
         c_default_data => "0",
         c_reg_last_bit => 1,
         c_addr_width => 0
      )
      PORT MAP (
         CLK => BU1729_CLK,
         D => BU1729_D,
         Q => BU1729_Q
      );

   BU1734_clk <= n152;
   BU1734_a(13) <= n574;
   BU1734_a(12) <= n575;
   BU1734_a(11) <= n576;
   BU1734_a(10) <= n577;
   BU1734_a(9) <= n578;
   BU1734_a(8) <= n579;
   BU1734_a(7) <= n580;
   BU1734_a(6) <= n581;
   BU1734_a(5) <= n582;
   BU1734_a(4) <= n583;
   BU1734_a(3) <= n584;
   BU1734_a(2) <= n585;
   BU1734_a(1) <= n586;
   BU1734_a(0) <= n587;
   BU1734_b(14) <= n616;
   BU1734_b(13) <= n617;
   BU1734_b(12) <= n618;
   BU1734_b(11) <= n619;
   BU1734_b(10) <= n620;
   BU1734_b(9) <= n621;
   BU1734_b(8) <= n622;
   BU1734_b(7) <= n623;
   BU1734_b(6) <= n624;
   BU1734_b(5) <= n625;
   BU1734_b(4) <= n626;
   BU1734_b(3) <= n627;
   BU1734_b(2) <= n628;
   BU1734_b(1) <= n629;
   BU1734_b(0) <= n630;
   n661 <= BU1734_q(28);
   n662 <= BU1734_q(27);
   n663 <= BU1734_q(26);
   n664 <= BU1734_q(25);
   n665 <= BU1734_q(24);
   n666 <= BU1734_q(23);
   n667 <= BU1734_q(22);
   n668 <= BU1734_q(21);
   n669 <= BU1734_q(20);
   n670 <= BU1734_q(19);
   n671 <= BU1734_q(18);
   n672 <= BU1734_q(17);
   n673 <= BU1734_q(16);
   n674 <= BU1734_q(15);
   n675 <= BU1734_q(14);
   n676 <= BU1734_q(13);
   n677 <= BU1734_q(12);
   n678 <= BU1734_q(11);
   n679 <= BU1734_q(10);
   n680 <= BU1734_q(9);
   n681 <= BU1734_q(8);
   n682 <= BU1734_q(7);
   n683 <= BU1734_q(6);
   n684 <= BU1734_q(5);
   n685 <= BU1734_q(4);
   n686 <= BU1734_q(3);
   n687 <= BU1734_q(2);
   n688 <= BU1734_q(1);
   n689 <= BU1734_q(0);
   BU1734_a_signed <= '0';
   BU1734_loadb <= '0';
   BU1734_swapb <= '0';
   BU1734_ce <= '1';
   BU1734_aclr <= '0';
   BU1734_sclr <= '0';
   BU1734_nd <= n338;
   BU1734 : mult_gen_v5_0
      GENERIC MAP (
         c_a_width => 14,
         c_out_width => 29,
         c_b_type => 0,
         c_has_b => 1,
         c_has_rdy => 1,
         bram_addr_width => 8,
         c_has_sclr => 0,
         c_has_nd => 1,
         c_reg_a_b_inputs => 1,
         c_enable_rlocs => 0,
         c_has_rfd => 1,
         c_mult_type => 1,
         c_has_swapb => 0,
         c_baat => 14,
         c_use_luts => 1,
         c_has_load_done => 0,
         c_has_a_signed => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 1,
         c_output_hold => 0,
         c_stack_adders => 0,
         c_mem_type => 0,
         c_b_constant => 0,
         c_has_q => 1,
         c_has_loadb => 0,
         c_pipeline => 1,
         c_has_o => 0,
         c_standalone => 1,
         c_mem_init_prefix => "mem",
         c_a_type => 0,
         c_b_width => 15,
         c_sqm_type => 0,
         c_b_value => "0"
      )
      PORT MAP (
         clk => BU1734_clk,
         a => BU1734_a,
         b => BU1734_b,
         o => BU1734_o,
         q => BU1734_q,
         a_signed => BU1734_a_signed,
         loadb => BU1734_loadb,
         load_done => BU1734_load_done,
         swapb => BU1734_swapb,
         ce => BU1734_ce,
         aclr => BU1734_aclr,
         sclr => BU1734_sclr,
         rfd => BU1734_rfd,
         nd => BU1734_nd,
         rdy => BU1734_rdy
      );

   BU1955_I(0) <= n689;
   BU1955_I(1) <= n688;
   BU1955_I(2) <= n687;
   BU1955_I(3) <= n686;
   BU1955_I(4) <= n685;
   n2187 <= BU1955_O;
   BU1955 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 5,
         c_input_inv_mask => "01111"
      )
      PORT MAP (
         I => BU1955_I,
         O => BU1955_O
      );

   BU1964_I0 <= n684;
   BU1964_I1 <= n685;
   BU1964_I2 <= n2187;
   BU1964_I3 <= '0';
   n2184 <= BU1964_O;
   BU1964 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU1964_I0,
         I1 => BU1964_I1,
         I2 => BU1964_I2,
         I3 => BU1964_I3,
         O => BU1964_O
      );

   BU1965_A(0) <= n684;
   BU1965_A(1) <= n683;
   BU1965_A(2) <= n682;
   BU1965_A(3) <= n681;
   BU1965_A(4) <= n680;
   BU1965_A(5) <= n679;
   BU1965_A(6) <= n678;
   BU1965_A(7) <= n677;
   BU1965_A(8) <= n676;
   BU1965_A(9) <= n675;
   BU1965_A(10) <= n674;
   BU1965_A(11) <= n673;
   BU1965_A(12) <= n672;
   BU1965_A(13) <= n671;
   BU1965_A(14) <= n670;
   BU1965_A(15) <= n669;
   BU1965_A(16) <= n668;
   BU1965_A(17) <= n667;
   BU1965_A(18) <= n666;
   BU1965_A(19) <= n665;
   BU1965_A(20) <= n664;
   BU1965_A(21) <= n663;
   BU1965_A(22) <= n662;
   BU1965_A(23) <= n661;
   BU1965_B(0) <= n2184;
   n2159 <= BU1965_S(0);
   n2160 <= BU1965_S(1);
   n2161 <= BU1965_S(2);
   n2162 <= BU1965_S(3);
   n2163 <= BU1965_S(4);
   n2164 <= BU1965_S(5);
   n2165 <= BU1965_S(6);
   n2166 <= BU1965_S(7);
   n2167 <= BU1965_S(8);
   n2168 <= BU1965_S(9);
   n2169 <= BU1965_S(10);
   n2170 <= BU1965_S(11);
   n2171 <= BU1965_S(12);
   n2172 <= BU1965_S(13);
   n2173 <= BU1965_S(14);
   n2174 <= BU1965_S(15);
   n2175 <= BU1965_S(16);
   n2176 <= BU1965_S(17);
   n2177 <= BU1965_S(18);
   n2178 <= BU1965_S(19);
   n2179 <= BU1965_S(20);
   n2180 <= BU1965_S(21);
   n2181 <= BU1965_S(22);
   n2182 <= BU1965_S(23);
   BU1965 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU1965_A,
         B => BU1965_B,
         S => BU1965_S
      );

   BU2066_I0 <= n661;
   BU2066_I1 <= n662;
   BU2066_I2 <= n2182;
   BU2066_I3 <= '0';
   n2193 <= BU2066_O;
   BU2066 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU2066_I0,
         I1 => BU2066_I1,
         I2 => BU2066_I2,
         I3 => BU2066_I3,
         O => BU2066_O
      );

   BU2068_I0 <= n661;
   BU2068_I1 <= n2182;
   BU2068_I2 <= '0';
   BU2068_I3 <= '0';
   n2195 <= BU2068_O;
   BU2068 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU2068_I0,
         I1 => BU2068_I1,
         I2 => BU2068_I2,
         I3 => BU2068_I3,
         O => BU2068_O
      );

   BU2069_D(0) <= n2159;
   BU2069_D(1) <= n2160;
   BU2069_D(2) <= n2161;
   BU2069_D(3) <= n2162;
   BU2069_D(4) <= n2163;
   BU2069_D(5) <= n2164;
   BU2069_D(6) <= n2165;
   BU2069_D(7) <= n2166;
   BU2069_D(8) <= n2167;
   BU2069_D(9) <= n2168;
   BU2069_D(10) <= n2169;
   BU2069_D(11) <= n2170;
   BU2069_D(12) <= n2171;
   BU2069_D(13) <= n2172;
   BU2069_D(14) <= n2173;
   BU2069_D(15) <= n2174;
   BU2069_D(16) <= n2175;
   BU2069_D(17) <= n2176;
   BU2069_D(18) <= n2177;
   BU2069_D(19) <= n2178;
   BU2069_D(20) <= n2179;
   BU2069_D(21) <= n2180;
   BU2069_D(22) <= n2181;
   n27 <= BU2069_Q(0);
   n28 <= BU2069_Q(1);
   n29 <= BU2069_Q(2);
   n30 <= BU2069_Q(3);
   n31 <= BU2069_Q(4);
   n32 <= BU2069_Q(5);
   n33 <= BU2069_Q(6);
   n34 <= BU2069_Q(7);
   n35 <= BU2069_Q(8);
   n36 <= BU2069_Q(9);
   n37 <= BU2069_Q(10);
   n38 <= BU2069_Q(11);
   n39 <= BU2069_Q(12);
   n40 <= BU2069_Q(13);
   n41 <= BU2069_Q(14);
   n42 <= BU2069_Q(15);
   n43 <= BU2069_Q(16);
   n44 <= BU2069_Q(17);
   n45 <= BU2069_Q(18);
   n46 <= BU2069_Q(19);
   n47 <= BU2069_Q(20);
   n48 <= BU2069_Q(21);
   n49 <= BU2069_Q(22);
   BU2069_CLK <= n152;
   BU2069_SCLR <= n2193;
   BU2069_SSET <= n2195;
   BU2069 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2069_D,
         Q => BU2069_Q,
         CLK => BU2069_CLK,
         SCLR => BU2069_SCLR,
         SSET => BU2069_SSET
      );

   BU2162_D(0) <= n2182;
   n50 <= BU2162_Q(0);
   BU2162_CLK <= n152;
   BU2162_SCLR <= n2195;
   BU2162_SSET <= n2193;
   BU2162 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2162_D,
         Q => BU2162_Q,
         CLK => BU2162_CLK,
         SCLR => BU2162_SCLR,
         SSET => BU2162_SSET
      );

   BU2457_D <= n2716;
   BU2457_C <= n152;
   BU2457_CE <= '1';
   n2674 <= BU2457_Q;
   BU2457 : FDE
      PORT MAP (
         D => BU2457_D,
         C => BU2457_C,
         CE => BU2457_CE,
         Q => BU2457_Q
      );

   BU2461_I(0) <= n2676;
   BU2461_I(1) <= n2677;
   BU2461_I(2) <= n2678;
   BU2461_I(3) <= n2679;
   BU2461_I(4) <= n2680;
   BU2461_I(5) <= n2681;
   BU2461_I(6) <= n2682;
   BU2461_I(7) <= n2683;
   BU2461_I(8) <= n2684;
   BU2461_I(9) <= n2685;
   BU2461_I(10) <= n2686;
   BU2461_I(11) <= n2687;
   BU2461_I(12) <= n2688;
   BU2461_I(13) <= n2689;
   BU2461_I(14) <= n2690;
   BU2461_I(15) <= n2691;
   n2943 <= BU2461_O;
   BU2461 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 16,
         c_input_inv_mask => "0111111111111111"
      )
      PORT MAP (
         I => BU2461_I,
         O => BU2461_O
      );

   BU2479_I0 <= n2692;
   BU2479_I1 <= n2691;
   BU2479_I2 <= n2943;
   BU2479_I3 <= '0';
   n2940 <= BU2479_O;
   BU2479 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU2479_I0,
         I1 => BU2479_I1,
         I2 => BU2479_I2,
         I3 => BU2479_I3,
         O => BU2479_O
      );

   BU2480_A(0) <= n2692;
   BU2480_A(1) <= n2693;
   BU2480_A(2) <= n2694;
   BU2480_A(3) <= n2695;
   BU2480_A(4) <= n2696;
   BU2480_A(5) <= n2697;
   BU2480_A(6) <= n2698;
   BU2480_A(7) <= n2699;
   BU2480_A(8) <= n2700;
   BU2480_A(9) <= n2701;
   BU2480_A(10) <= n2702;
   BU2480_A(11) <= n2703;
   BU2480_A(12) <= n2704;
   BU2480_A(13) <= n2705;
   BU2480_A(14) <= n2706;
   BU2480_A(15) <= n2707;
   BU2480_A(16) <= n2708;
   BU2480_A(17) <= n2709;
   BU2480_A(18) <= n2710;
   BU2480_A(19) <= n2711;
   BU2480_A(20) <= n2712;
   BU2480_A(21) <= n2713;
   BU2480_A(22) <= n2714;
   BU2480_A(23) <= n2715;
   BU2480_B(0) <= n2940;
   n2915 <= BU2480_S(0);
   n2916 <= BU2480_S(1);
   n2917 <= BU2480_S(2);
   n2918 <= BU2480_S(3);
   n2919 <= BU2480_S(4);
   n2920 <= BU2480_S(5);
   n2921 <= BU2480_S(6);
   n2922 <= BU2480_S(7);
   n2923 <= BU2480_S(8);
   n2924 <= BU2480_S(9);
   n2925 <= BU2480_S(10);
   n2926 <= BU2480_S(11);
   n2927 <= BU2480_S(12);
   n2928 <= BU2480_S(13);
   n2929 <= BU2480_S(14);
   n2930 <= BU2480_S(15);
   n2931 <= BU2480_S(16);
   n2932 <= BU2480_S(17);
   n2933 <= BU2480_S(18);
   n2934 <= BU2480_S(19);
   n2935 <= BU2480_S(20);
   n2936 <= BU2480_S(21);
   n2937 <= BU2480_S(22);
   n2938 <= BU2480_S(23);
   BU2480 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU2480_A,
         B => BU2480_B,
         S => BU2480_S
      );

   BU2581_I0 <= n2715;
   BU2581_I1 <= n2714;
   BU2581_I2 <= n2938;
   BU2581_I3 <= '0';
   n2960 <= BU2581_O;
   BU2581 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU2581_I0,
         I1 => BU2581_I1,
         I2 => BU2581_I2,
         I3 => BU2581_I3,
         O => BU2581_O
      );

   BU2583_I0 <= n2715;
   BU2583_I1 <= n2938;
   BU2583_I2 <= '0';
   BU2583_I3 <= '0';
   n2962 <= BU2583_O;
   BU2583 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU2583_I0,
         I1 => BU2583_I1,
         I2 => BU2583_I2,
         I3 => BU2583_I3,
         O => BU2583_O
      );

   BU2584_D(0) <= n2915;
   BU2584_D(1) <= n2916;
   BU2584_D(2) <= n2917;
   BU2584_D(3) <= n2918;
   BU2584_D(4) <= n2919;
   BU2584_D(5) <= n2920;
   BU2584_D(6) <= n2921;
   BU2584_D(7) <= n2922;
   BU2584_D(8) <= n2923;
   BU2584_D(9) <= n2924;
   BU2584_D(10) <= n2925;
   BU2584_D(11) <= n2926;
   BU2584_D(12) <= n2927;
   BU2584_D(13) <= n2928;
   BU2584_D(14) <= n2929;
   BU2584_D(15) <= n2930;
   BU2584_D(16) <= n2931;
   BU2584_D(17) <= n2932;
   BU2584_D(18) <= n2933;
   BU2584_D(19) <= n2934;
   BU2584_D(20) <= n2935;
   BU2584_D(21) <= n2936;
   BU2584_D(22) <= n2937;
   n2602 <= BU2584_Q(0);
   n2603 <= BU2584_Q(1);
   n2604 <= BU2584_Q(2);
   n2605 <= BU2584_Q(3);
   n2606 <= BU2584_Q(4);
   n2607 <= BU2584_Q(5);
   n2608 <= BU2584_Q(6);
   n2609 <= BU2584_Q(7);
   n2610 <= BU2584_Q(8);
   n2611 <= BU2584_Q(9);
   n2612 <= BU2584_Q(10);
   n2613 <= BU2584_Q(11);
   n2614 <= BU2584_Q(12);
   n2615 <= BU2584_Q(13);
   n2616 <= BU2584_Q(14);
   n2617 <= BU2584_Q(15);
   n2618 <= BU2584_Q(16);
   n2619 <= BU2584_Q(17);
   n2620 <= BU2584_Q(18);
   n2621 <= BU2584_Q(19);
   n2622 <= BU2584_Q(20);
   n2623 <= BU2584_Q(21);
   n2624 <= BU2584_Q(22);
   BU2584_CLK <= n152;
   BU2584_SCLR <= n2960;
   BU2584_SSET <= n2962;
   BU2584 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2584_D,
         Q => BU2584_Q,
         CLK => BU2584_CLK,
         SCLR => BU2584_SCLR,
         SSET => BU2584_SSET
      );

   BU2677_D(0) <= n2938;
   n2625 <= BU2677_Q(0);
   BU2677_CLK <= n152;
   BU2677_SCLR <= n2962;
   BU2677_SSET <= n2960;
   BU2677 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU2677_D,
         Q => BU2677_Q,
         CLK => BU2677_CLK,
         SCLR => BU2677_SCLR,
         SSET => BU2677_SSET
      );

   BU6771_I(0) <= n2717;
   BU6771_I(1) <= n2718;
   BU6771_I(2) <= n2719;
   BU6771_I(3) <= n2720;
   BU6771_I(4) <= n2721;
   BU6771_I(5) <= n2722;
   BU6771_I(6) <= n2723;
   BU6771_I(7) <= n2724;
   BU6771_I(8) <= n2725;
   BU6771_I(9) <= n2726;
   BU6771_I(10) <= n2727;
   BU6771_I(11) <= n2728;
   BU6771_I(12) <= n2729;
   BU6771_I(13) <= n2730;
   BU6771_I(14) <= n2731;
   BU6771_I(15) <= n2732;
   n3431 <= BU6771_O;
   BU6771 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 16,
         c_input_inv_mask => "0111111111111111"
      )
      PORT MAP (
         I => BU6771_I,
         O => BU6771_O
      );

   BU6789_I0 <= n2733;
   BU6789_I1 <= n2732;
   BU6789_I2 <= n3431;
   BU6789_I3 <= '0';
   n3428 <= BU6789_O;
   BU6789 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU6789_I0,
         I1 => BU6789_I1,
         I2 => BU6789_I2,
         I3 => BU6789_I3,
         O => BU6789_O
      );

   BU6790_A(0) <= n2733;
   BU6790_A(1) <= n2734;
   BU6790_A(2) <= n2735;
   BU6790_A(3) <= n2736;
   BU6790_A(4) <= n2737;
   BU6790_A(5) <= n2738;
   BU6790_A(6) <= n2739;
   BU6790_A(7) <= n2740;
   BU6790_A(8) <= n2741;
   BU6790_A(9) <= n2742;
   BU6790_A(10) <= n2743;
   BU6790_A(11) <= n2744;
   BU6790_A(12) <= n2745;
   BU6790_A(13) <= n2746;
   BU6790_A(14) <= n2747;
   BU6790_A(15) <= n2748;
   BU6790_A(16) <= n2749;
   BU6790_A(17) <= n2750;
   BU6790_A(18) <= n2751;
   BU6790_A(19) <= n2752;
   BU6790_A(20) <= n2753;
   BU6790_A(21) <= n2754;
   BU6790_A(22) <= n2755;
   BU6790_A(23) <= n2756;
   BU6790_B(0) <= n3428;
   n3403 <= BU6790_S(0);
   n3404 <= BU6790_S(1);
   n3405 <= BU6790_S(2);
   n3406 <= BU6790_S(3);
   n3407 <= BU6790_S(4);
   n3408 <= BU6790_S(5);
   n3409 <= BU6790_S(6);
   n3410 <= BU6790_S(7);
   n3411 <= BU6790_S(8);
   n3412 <= BU6790_S(9);
   n3413 <= BU6790_S(10);
   n3414 <= BU6790_S(11);
   n3415 <= BU6790_S(12);
   n3416 <= BU6790_S(13);
   n3417 <= BU6790_S(14);
   n3418 <= BU6790_S(15);
   n3419 <= BU6790_S(16);
   n3420 <= BU6790_S(17);
   n3421 <= BU6790_S(18);
   n3422 <= BU6790_S(19);
   n3423 <= BU6790_S(20);
   n3424 <= BU6790_S(21);
   n3425 <= BU6790_S(22);
   n3426 <= BU6790_S(23);
   BU6790 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 24,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 25,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 24,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU6790_A,
         B => BU6790_B,
         S => BU6790_S
      );

   BU6891_I0 <= n2756;
   BU6891_I1 <= n2755;
   BU6891_I2 <= n3426;
   BU6891_I3 <= '0';
   n3448 <= BU6891_O;
   BU6891 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU6891_I0,
         I1 => BU6891_I1,
         I2 => BU6891_I2,
         I3 => BU6891_I3,
         O => BU6891_O
      );

   BU6893_I0 <= n2756;
   BU6893_I1 <= n3426;
   BU6893_I2 <= '0';
   BU6893_I3 <= '0';
   n3450 <= BU6893_O;
   BU6893 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU6893_I0,
         I1 => BU6893_I1,
         I2 => BU6893_I2,
         I3 => BU6893_I3,
         O => BU6893_O
      );

   BU6894_D(0) <= n3403;
   BU6894_D(1) <= n3404;
   BU6894_D(2) <= n3405;
   BU6894_D(3) <= n3406;
   BU6894_D(4) <= n3407;
   BU6894_D(5) <= n3408;
   BU6894_D(6) <= n3409;
   BU6894_D(7) <= n3410;
   BU6894_D(8) <= n3411;
   BU6894_D(9) <= n3412;
   BU6894_D(10) <= n3413;
   BU6894_D(11) <= n3414;
   BU6894_D(12) <= n3415;
   BU6894_D(13) <= n3416;
   BU6894_D(14) <= n3417;
   BU6894_D(15) <= n3418;
   BU6894_D(16) <= n3419;
   BU6894_D(17) <= n3420;
   BU6894_D(18) <= n3421;
   BU6894_D(19) <= n3422;
   BU6894_D(20) <= n3423;
   BU6894_D(21) <= n3424;
   BU6894_D(22) <= n3425;
   n2626 <= BU6894_Q(0);
   n2627 <= BU6894_Q(1);
   n2628 <= BU6894_Q(2);
   n2629 <= BU6894_Q(3);
   n2630 <= BU6894_Q(4);
   n2631 <= BU6894_Q(5);
   n2632 <= BU6894_Q(6);
   n2633 <= BU6894_Q(7);
   n2634 <= BU6894_Q(8);
   n2635 <= BU6894_Q(9);
   n2636 <= BU6894_Q(10);
   n2637 <= BU6894_Q(11);
   n2638 <= BU6894_Q(12);
   n2639 <= BU6894_Q(13);
   n2640 <= BU6894_Q(14);
   n2641 <= BU6894_Q(15);
   n2642 <= BU6894_Q(16);
   n2643 <= BU6894_Q(17);
   n2644 <= BU6894_Q(18);
   n2645 <= BU6894_Q(19);
   n2646 <= BU6894_Q(20);
   n2647 <= BU6894_Q(21);
   n2648 <= BU6894_Q(22);
   BU6894_CLK <= n152;
   BU6894_SCLR <= n3448;
   BU6894_SSET <= n3450;
   BU6894 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 23,
         c_has_ce => 0,
         c_sinit_val => "00000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU6894_D,
         Q => BU6894_Q,
         CLK => BU6894_CLK,
         SCLR => BU6894_SCLR,
         SSET => BU6894_SSET
      );

   BU6987_D(0) <= n3426;
   n2649 <= BU6987_Q(0);
   BU6987_CLK <= n152;
   BU6987_SCLR <= n3450;
   BU6987_SSET <= n3448;
   BU6987 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU6987_D,
         Q => BU6987_Q,
         CLK => BU6987_CLK,
         SCLR => BU6987_SCLR,
         SSET => BU6987_SSET
      );

   BU2173_D <= n2626;
   BU2173_C <= n152;
   BU2173_CE <= '1';
   n2650 <= BU2173_Q;
   BU2173 : FDE
      PORT MAP (
         D => BU2173_D,
         C => BU2173_C,
         CE => BU2173_CE,
         Q => BU2173_Q
      );

   BU2175_D <= n2627;
   BU2175_C <= n152;
   BU2175_CE <= '1';
   n2651 <= BU2175_Q;
   BU2175 : FDE
      PORT MAP (
         D => BU2175_D,
         C => BU2175_C,
         CE => BU2175_CE,
         Q => BU2175_Q
      );

   BU2177_D <= n2628;
   BU2177_C <= n152;
   BU2177_CE <= '1';
   n2652 <= BU2177_Q;
   BU2177 : FDE
      PORT MAP (
         D => BU2177_D,
         C => BU2177_C,
         CE => BU2177_CE,
         Q => BU2177_Q
      );

   BU2179_D <= n2629;
   BU2179_C <= n152;
   BU2179_CE <= '1';
   n2653 <= BU2179_Q;
   BU2179 : FDE
      PORT MAP (
         D => BU2179_D,
         C => BU2179_C,
         CE => BU2179_CE,
         Q => BU2179_Q
      );

   BU2181_D <= n2630;
   BU2181_C <= n152;
   BU2181_CE <= '1';
   n2654 <= BU2181_Q;
   BU2181 : FDE
      PORT MAP (
         D => BU2181_D,
         C => BU2181_C,
         CE => BU2181_CE,
         Q => BU2181_Q
      );

   BU2183_D <= n2631;
   BU2183_C <= n152;
   BU2183_CE <= '1';
   n2655 <= BU2183_Q;
   BU2183 : FDE
      PORT MAP (
         D => BU2183_D,
         C => BU2183_C,
         CE => BU2183_CE,
         Q => BU2183_Q
      );

   BU2185_D <= n2632;
   BU2185_C <= n152;
   BU2185_CE <= '1';
   n2656 <= BU2185_Q;
   BU2185 : FDE
      PORT MAP (
         D => BU2185_D,
         C => BU2185_C,
         CE => BU2185_CE,
         Q => BU2185_Q
      );

   BU2187_D <= n2633;
   BU2187_C <= n152;
   BU2187_CE <= '1';
   n2657 <= BU2187_Q;
   BU2187 : FDE
      PORT MAP (
         D => BU2187_D,
         C => BU2187_C,
         CE => BU2187_CE,
         Q => BU2187_Q
      );

   BU2189_D <= n2634;
   BU2189_C <= n152;
   BU2189_CE <= '1';
   n2658 <= BU2189_Q;
   BU2189 : FDE
      PORT MAP (
         D => BU2189_D,
         C => BU2189_C,
         CE => BU2189_CE,
         Q => BU2189_Q
      );

   BU2191_D <= n2635;
   BU2191_C <= n152;
   BU2191_CE <= '1';
   n2659 <= BU2191_Q;
   BU2191 : FDE
      PORT MAP (
         D => BU2191_D,
         C => BU2191_C,
         CE => BU2191_CE,
         Q => BU2191_Q
      );

   BU2193_D <= n2636;
   BU2193_C <= n152;
   BU2193_CE <= '1';
   n2660 <= BU2193_Q;
   BU2193 : FDE
      PORT MAP (
         D => BU2193_D,
         C => BU2193_C,
         CE => BU2193_CE,
         Q => BU2193_Q
      );

   BU2195_D <= n2637;
   BU2195_C <= n152;
   BU2195_CE <= '1';
   n2661 <= BU2195_Q;
   BU2195 : FDE
      PORT MAP (
         D => BU2195_D,
         C => BU2195_C,
         CE => BU2195_CE,
         Q => BU2195_Q
      );

   BU2197_D <= n2638;
   BU2197_C <= n152;
   BU2197_CE <= '1';
   n2662 <= BU2197_Q;
   BU2197 : FDE
      PORT MAP (
         D => BU2197_D,
         C => BU2197_C,
         CE => BU2197_CE,
         Q => BU2197_Q
      );

   BU2199_D <= n2639;
   BU2199_C <= n152;
   BU2199_CE <= '1';
   n2663 <= BU2199_Q;
   BU2199 : FDE
      PORT MAP (
         D => BU2199_D,
         C => BU2199_C,
         CE => BU2199_CE,
         Q => BU2199_Q
      );

   BU2201_D <= n2640;
   BU2201_C <= n152;
   BU2201_CE <= '1';
   n2664 <= BU2201_Q;
   BU2201 : FDE
      PORT MAP (
         D => BU2201_D,
         C => BU2201_C,
         CE => BU2201_CE,
         Q => BU2201_Q
      );

   BU2203_D <= n2641;
   BU2203_C <= n152;
   BU2203_CE <= '1';
   n2665 <= BU2203_Q;
   BU2203 : FDE
      PORT MAP (
         D => BU2203_D,
         C => BU2203_C,
         CE => BU2203_CE,
         Q => BU2203_Q
      );

   BU2205_D <= n2642;
   BU2205_C <= n152;
   BU2205_CE <= '1';
   n2666 <= BU2205_Q;
   BU2205 : FDE
      PORT MAP (
         D => BU2205_D,
         C => BU2205_C,
         CE => BU2205_CE,
         Q => BU2205_Q
      );

   BU2207_D <= n2643;
   BU2207_C <= n152;
   BU2207_CE <= '1';
   n2667 <= BU2207_Q;
   BU2207 : FDE
      PORT MAP (
         D => BU2207_D,
         C => BU2207_C,
         CE => BU2207_CE,
         Q => BU2207_Q
      );

   BU2209_D <= n2644;
   BU2209_C <= n152;
   BU2209_CE <= '1';
   n2668 <= BU2209_Q;
   BU2209 : FDE
      PORT MAP (
         D => BU2209_D,
         C => BU2209_C,
         CE => BU2209_CE,
         Q => BU2209_Q
      );

   BU2211_D <= n2645;
   BU2211_C <= n152;
   BU2211_CE <= '1';
   n2669 <= BU2211_Q;
   BU2211 : FDE
      PORT MAP (
         D => BU2211_D,
         C => BU2211_C,
         CE => BU2211_CE,
         Q => BU2211_Q
      );

   BU2213_D <= n2646;
   BU2213_C <= n152;
   BU2213_CE <= '1';
   n2670 <= BU2213_Q;
   BU2213 : FDE
      PORT MAP (
         D => BU2213_D,
         C => BU2213_C,
         CE => BU2213_CE,
         Q => BU2213_Q
      );

   BU2215_D <= n2647;
   BU2215_C <= n152;
   BU2215_CE <= '1';
   n2671 <= BU2215_Q;
   BU2215 : FDE
      PORT MAP (
         D => BU2215_D,
         C => BU2215_C,
         CE => BU2215_CE,
         Q => BU2215_Q
      );

   BU2217_D <= n2648;
   BU2217_C <= n152;
   BU2217_CE <= '1';
   n2672 <= BU2217_Q;
   BU2217 : FDE
      PORT MAP (
         D => BU2217_D,
         C => BU2217_C,
         CE => BU2217_CE,
         Q => BU2217_Q
      );

   BU2219_D <= n2649;
   BU2219_C <= n152;
   BU2219_CE <= '1';
   n2673 <= BU2219_Q;
   BU2219 : FDE
      PORT MAP (
         D => BU2219_D,
         C => BU2219_C,
         CE => BU2219_CE,
         Q => BU2219_Q
      );

   BU2220_MA(0) <= n2650;
   BU2220_MA(1) <= n2651;
   BU2220_MA(2) <= n2652;
   BU2220_MA(3) <= n2653;
   BU2220_MA(4) <= n2654;
   BU2220_MA(5) <= n2655;
   BU2220_MA(6) <= n2656;
   BU2220_MA(7) <= n2657;
   BU2220_MA(8) <= n2658;
   BU2220_MA(9) <= n2659;
   BU2220_MA(10) <= n2660;
   BU2220_MA(11) <= n2661;
   BU2220_MA(12) <= n2662;
   BU2220_MA(13) <= n2663;
   BU2220_MA(14) <= n2664;
   BU2220_MA(15) <= n2665;
   BU2220_MA(16) <= n2666;
   BU2220_MA(17) <= n2667;
   BU2220_MA(18) <= n2668;
   BU2220_MA(19) <= n2669;
   BU2220_MA(20) <= n2670;
   BU2220_MA(21) <= n2671;
   BU2220_MA(22) <= n2672;
   BU2220_MA(23) <= n2673;
   BU2220_MB(0) <= n2602;
   BU2220_MB(1) <= n2603;
   BU2220_MB(2) <= n2604;
   BU2220_MB(3) <= n2605;
   BU2220_MB(4) <= n2606;
   BU2220_MB(5) <= n2607;
   BU2220_MB(6) <= n2608;
   BU2220_MB(7) <= n2609;
   BU2220_MB(8) <= n2610;
   BU2220_MB(9) <= n2611;
   BU2220_MB(10) <= n2612;
   BU2220_MB(11) <= n2613;
   BU2220_MB(12) <= n2614;
   BU2220_MB(13) <= n2615;
   BU2220_MB(14) <= n2616;
   BU2220_MB(15) <= n2617;
   BU2220_MB(16) <= n2618;
   BU2220_MB(17) <= n2619;
   BU2220_MB(18) <= n2620;
   BU2220_MB(19) <= n2621;
   BU2220_MB(20) <= n2622;
   BU2220_MB(21) <= n2623;
   BU2220_MB(22) <= n2624;
   BU2220_MB(23) <= n2625;
   BU2220_S(0) <= n2674;
   n56 <= BU2220_Q(0);
   n57 <= BU2220_Q(1);
   n58 <= BU2220_Q(2);
   n59 <= BU2220_Q(3);
   n60 <= BU2220_Q(4);
   n61 <= BU2220_Q(5);
   n62 <= BU2220_Q(6);
   n63 <= BU2220_Q(7);
   n64 <= BU2220_Q(8);
   n65 <= BU2220_Q(9);
   n66 <= BU2220_Q(10);
   n67 <= BU2220_Q(11);
   n68 <= BU2220_Q(12);
   n69 <= BU2220_Q(13);
   n70 <= BU2220_Q(14);
   n71 <= BU2220_Q(15);
   n72 <= BU2220_Q(16);
   n73 <= BU2220_Q(17);
   n74 <= BU2220_Q(18);
   n75 <= BU2220_Q(19);
   n76 <= BU2220_Q(20);
   n77 <= BU2220_Q(21);
   n78 <= BU2220_Q(22);
   n79 <= BU2220_Q(23);
   BU2220_CLK <= n152;
   BU2220 : C_MUX_BUS_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_has_en => 0,
         c_sync_priority => 0,
         c_has_sclr => 0,
         c_width => 24,
         c_enable_rlocs => 0,
         c_sel_width => 1,
         c_latency => 1,
         c_ainit_val => "000000000000000000000000",
         c_has_ce => 0,
         c_mux_type => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "000000000000000000000000",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 1,
         c_has_o => 0,
         c_inputs => 2
      )
      PORT MAP (
         MA => BU2220_MA,
         MB => BU2220_MB,
         S => BU2220_S,
         Q => BU2220_Q,
         CLK => BU2220_CLK
      );

   BU2448_D <= n2674;
   BU2448_C <= n152;
   BU2448_CE <= '1';
   n2675 <= BU2448_Q;
   BU2448 : FDE
      PORT MAP (
         D => BU2448_D,
         C => BU2448_C,
         CE => BU2448_CE,
         Q => BU2448_Q
      );

   BU2452_I0 <= n2674;
   BU2452_I1 <= n2675;
   BU2452_I2 <= '0';
   BU2452_I3 <= '0';
   n4288 <= BU2452_O;
   BU2452 : LUT4
      GENERIC MAP (
         INIT  => X"eeee"
      )
      PORT MAP (
         I0 => BU2452_I0,
         I1 => BU2452_I1,
         I2 => BU2452_I2,
         I3 => BU2452_I3,
         O => BU2452_O
      );

   BU2453_D <= n4288;
   BU2453_C <= n152;
   BU2453_CE <= '1';
   n55 <= BU2453_Q;
   BU2453 : FDE
      PORT MAP (
         D => BU2453_D,
         C => BU2453_C,
         CE => BU2453_CE,
         Q => BU2453_Q
      );

   BU2682_DIN(0) <= n3;
   BU2682_DIN(1) <= n4;
   BU2682_DIN(2) <= n5;
   BU2682_DIN(3) <= n6;
   BU2682_DIN(4) <= n7;
   BU2682_DIN(5) <= n8;
   BU2682_DIN(6) <= n9;
   BU2682_DIN(7) <= n10;
   BU2682_DIN(8) <= n11;
   BU2682_DIN(9) <= n12;
   BU2682_DIN(10) <= n13;
   BU2682_DIN(11) <= n14;
   BU2682_DIN(12) <= n15;
   BU2682_DIN(13) <= n16;
   BU2682_DIN(14) <= n17;
   BU2682_DIN(15) <= n18;
   BU2682_DIN(16) <= n19;
   BU2682_DIN(17) <= n20;
   BU2682_DIN(18) <= n21;
   BU2682_DIN(19) <= n22;
   BU2682_DIN(20) <= n23;
   BU2682_DIN(21) <= n24;
   BU2682_DIN(22) <= n25;
   BU2682_DIN(23) <= n26;
   BU2682_ND <= n2;
   BU2682_CLK <= n152;
   n2676 <= BU2682_DOUT(0);
   n2677 <= BU2682_DOUT(1);
   n2678 <= BU2682_DOUT(2);
   n2679 <= BU2682_DOUT(3);
   n2680 <= BU2682_DOUT(4);
   n2681 <= BU2682_DOUT(5);
   n2682 <= BU2682_DOUT(6);
   n2683 <= BU2682_DOUT(7);
   n2684 <= BU2682_DOUT(8);
   n2685 <= BU2682_DOUT(9);
   n2686 <= BU2682_DOUT(10);
   n2687 <= BU2682_DOUT(11);
   n2688 <= BU2682_DOUT(12);
   n2689 <= BU2682_DOUT(13);
   n2690 <= BU2682_DOUT(14);
   n2691 <= BU2682_DOUT(15);
   n2692 <= BU2682_DOUT(16);
   n2693 <= BU2682_DOUT(17);
   n2694 <= BU2682_DOUT(18);
   n2695 <= BU2682_DOUT(19);
   n2696 <= BU2682_DOUT(20);
   n2697 <= BU2682_DOUT(21);
   n2698 <= BU2682_DOUT(22);
   n2699 <= BU2682_DOUT(23);
   n2700 <= BU2682_DOUT(24);
   n2701 <= BU2682_DOUT(25);
   n2702 <= BU2682_DOUT(26);
   n2703 <= BU2682_DOUT(27);
   n2704 <= BU2682_DOUT(28);
   n2705 <= BU2682_DOUT(29);
   n2706 <= BU2682_DOUT(30);
   n2707 <= BU2682_DOUT(31);
   n2708 <= BU2682_DOUT(32);
   n2709 <= BU2682_DOUT(33);
   n2710 <= BU2682_DOUT(34);
   n2711 <= BU2682_DOUT(35);
   n2712 <= BU2682_DOUT(36);
   n2713 <= BU2682_DOUT(37);
   n2714 <= BU2682_DOUT(38);
   n2715 <= BU2682_DOUT(39);
   n2716 <= BU2682_RDY;
   BU2682 : C_CIC_V3_0
      GENERIC MAP (
         c_differential_delay => 1,
         c_sample_rate_change_max => 16383,
         c_number_channels => 1,
         c_filter_type => 2,
         c_result_width => 40,
         c_enable_rlocs => 0,
         c_sample_rate_change => 5,
         c_latency => 1,
         c_sample_rate_change_min => 4,
         c_sample_rate_change_type => 2,
         c_data_width => 24,
         c_stages => 7
      )
      PORT MAP (
         DIN => BU2682_DIN,
         ND => BU2682_ND,
         RFD => BU2682_RFD,
         CLK => BU2682_CLK,
         DOUT => BU2682_DOUT,
         RDY => BU2682_RDY
      );

   BU6992_DIN(0) <= n27;
   BU6992_DIN(1) <= n28;
   BU6992_DIN(2) <= n29;
   BU6992_DIN(3) <= n30;
   BU6992_DIN(4) <= n31;
   BU6992_DIN(5) <= n32;
   BU6992_DIN(6) <= n33;
   BU6992_DIN(7) <= n34;
   BU6992_DIN(8) <= n35;
   BU6992_DIN(9) <= n36;
   BU6992_DIN(10) <= n37;
   BU6992_DIN(11) <= n38;
   BU6992_DIN(12) <= n39;
   BU6992_DIN(13) <= n40;
   BU6992_DIN(14) <= n41;
   BU6992_DIN(15) <= n42;
   BU6992_DIN(16) <= n43;
   BU6992_DIN(17) <= n44;
   BU6992_DIN(18) <= n45;
   BU6992_DIN(19) <= n46;
   BU6992_DIN(20) <= n47;
   BU6992_DIN(21) <= n48;
   BU6992_DIN(22) <= n49;
   BU6992_DIN(23) <= n50;
   BU6992_ND <= n2;
   BU6992_CLK <= n152;
   n2717 <= BU6992_DOUT(0);
   n2718 <= BU6992_DOUT(1);
   n2719 <= BU6992_DOUT(2);
   n2720 <= BU6992_DOUT(3);
   n2721 <= BU6992_DOUT(4);
   n2722 <= BU6992_DOUT(5);
   n2723 <= BU6992_DOUT(6);
   n2724 <= BU6992_DOUT(7);
   n2725 <= BU6992_DOUT(8);
   n2726 <= BU6992_DOUT(9);
   n2727 <= BU6992_DOUT(10);
   n2728 <= BU6992_DOUT(11);
   n2729 <= BU6992_DOUT(12);
   n2730 <= BU6992_DOUT(13);
   n2731 <= BU6992_DOUT(14);
   n2732 <= BU6992_DOUT(15);
   n2733 <= BU6992_DOUT(16);
   n2734 <= BU6992_DOUT(17);
   n2735 <= BU6992_DOUT(18);
   n2736 <= BU6992_DOUT(19);
   n2737 <= BU6992_DOUT(20);
   n2738 <= BU6992_DOUT(21);
   n2739 <= BU6992_DOUT(22);
   n2740 <= BU6992_DOUT(23);
   n2741 <= BU6992_DOUT(24);
   n2742 <= BU6992_DOUT(25);
   n2743 <= BU6992_DOUT(26);
   n2744 <= BU6992_DOUT(27);
   n2745 <= BU6992_DOUT(28);
   n2746 <= BU6992_DOUT(29);
   n2747 <= BU6992_DOUT(30);
   n2748 <= BU6992_DOUT(31);
   n2749 <= BU6992_DOUT(32);
   n2750 <= BU6992_DOUT(33);
   n2751 <= BU6992_DOUT(34);
   n2752 <= BU6992_DOUT(35);
   n2753 <= BU6992_DOUT(36);
   n2754 <= BU6992_DOUT(37);
   n2755 <= BU6992_DOUT(38);
   n2756 <= BU6992_DOUT(39);
   BU6992 : C_CIC_V3_0
      GENERIC MAP (
         c_differential_delay => 1,
         c_sample_rate_change_max => 16383,
         c_number_channels => 1,
         c_filter_type => 2,
         c_result_width => 40,
         c_enable_rlocs => 0,
         c_sample_rate_change => 5,
         c_latency => 1,
         c_sample_rate_change_min => 4,
         c_sample_rate_change_type => 2,
         c_data_width => 24,
         c_stages => 7
      )
      PORT MAP (
         DIN => BU6992_DIN,
         ND => BU6992_ND,
         RFD => BU6992_RFD,
         CLK => BU6992_CLK,
         DOUT => BU6992_DOUT,
         RDY => BU6992_RDY
      );

   BU11080_ND <= n55;
   n6252 <= BU11080_RDY;
   BU11080_CLK <= n152;
   BU11080_DIN(0) <= n56;
   BU11080_DIN(1) <= n57;
   BU11080_DIN(2) <= n58;
   BU11080_DIN(3) <= n59;
   BU11080_DIN(4) <= n60;
   BU11080_DIN(5) <= n61;
   BU11080_DIN(6) <= n62;
   BU11080_DIN(7) <= n63;
   BU11080_DIN(8) <= n64;
   BU11080_DIN(9) <= n65;
   BU11080_DIN(10) <= n66;
   BU11080_DIN(11) <= n67;
   BU11080_DIN(12) <= n68;
   BU11080_DIN(13) <= n69;
   BU11080_DIN(14) <= n70;
   BU11080_DIN(15) <= n71;
   BU11080_DIN(16) <= n72;
   BU11080_DIN(17) <= n73;
   BU11080_DIN(18) <= n74;
   BU11080_DIN(19) <= n75;
   BU11080_DIN(20) <= n76;
   BU11080_DIN(21) <= n77;
   BU11080_DIN(22) <= n78;
   BU11080_DIN(23) <= n79;
   n6210 <= BU11080_DOUT(0);
   n6211 <= BU11080_DOUT(1);
   n6212 <= BU11080_DOUT(2);
   n6213 <= BU11080_DOUT(3);
   n6214 <= BU11080_DOUT(4);
   n6215 <= BU11080_DOUT(5);
   n6216 <= BU11080_DOUT(6);
   n6217 <= BU11080_DOUT(7);
   n6218 <= BU11080_DOUT(8);
   n6219 <= BU11080_DOUT(9);
   n6220 <= BU11080_DOUT(10);
   n6221 <= BU11080_DOUT(11);
   n6222 <= BU11080_DOUT(12);
   n6223 <= BU11080_DOUT(13);
   n6224 <= BU11080_DOUT(14);
   n6225 <= BU11080_DOUT(15);
   n6226 <= BU11080_DOUT(16);
   n6227 <= BU11080_DOUT(17);
   n6228 <= BU11080_DOUT(18);
   n6229 <= BU11080_DOUT(19);
   n6230 <= BU11080_DOUT(20);
   n6231 <= BU11080_DOUT(21);
   n6232 <= BU11080_DOUT(22);
   n6233 <= BU11080_DOUT(23);
   n6234 <= BU11080_DOUT(24);
   n6235 <= BU11080_DOUT(25);
   n6236 <= BU11080_DOUT(26);
   n6237 <= BU11080_DOUT(27);
   n6238 <= BU11080_DOUT(28);
   n6239 <= BU11080_DOUT(29);
   n6240 <= BU11080_DOUT(30);
   n6241 <= BU11080_DOUT(31);
   n6242 <= BU11080_DOUT(32);
   n6243 <= BU11080_DOUT(33);
   n6244 <= BU11080_DOUT(34);
   n6245 <= BU11080_DOUT(35);
   n6246 <= BU11080_DOUT(36);
   n6247 <= BU11080_DOUT(37);
   n6248 <= BU11080_DOUT(38);
   n6249 <= BU11080_DOUT(39);
   n6250 <= BU11080_DOUT(40);
   n6251 <= BU11080_DOUT(41);
   BU11080 : C_DA_FIR_V7_0
      GENERIC MAP (
         c_has_sout_r => 0,
         c_result_width => 42,
         c_reload_delay => 401,
         c_data_type => 0,
         c_filter_type => 2,
         c_channels => 2,
         c_response => 0,
         c_has_sout_f => 0,
         c_reg_output => 0,
         c_taps => 46,
         c_data_width => 24,
         c_enable_rlocs => 0,
         c_coeff_type => 0,
         c_reload_mem_type => 2,
         c_has_sin_r => 0,
         c_reload => 0,
         c_baat => 7,
         c_latency => 15,
         c_coeff_width => 16,
         c_optimize => 1,
         c_use_model_func => 0,
         c_zpf => 1,
         c_has_sin_f => 0,
         c_shape => 0,
         c_saturate => 0,
         c_has_sel_o => 0,
         c_mem_init_file => "ddcv1_0_CFIR.mif",
         c_polyphase_factor => 2,
         c_has_sel_i => 0,
         c_has_reset => 0
      )
      PORT MAP (
         ND => BU11080_ND,
         RDY => BU11080_RDY,
         CLK => BU11080_CLK,
         RFD => BU11080_RFD,
         DIN => BU11080_DIN,
         DOUT => BU11080_DOUT
      );

   BU20456_I(0) <= n6210;
   BU20456_I(1) <= n6211;
   BU20456_I(2) <= n6212;
   BU20456_I(3) <= n6213;
   BU20456_I(4) <= n6214;
   BU20456_I(5) <= n6215;
   BU20456_I(6) <= n6216;
   BU20456_I(7) <= n6217;
   BU20456_I(8) <= n6218;
   BU20456_I(9) <= n6219;
   BU20456_I(10) <= n6220;
   BU20456_I(11) <= n6221;
   BU20456_I(12) <= n6222;
   BU20456_I(13) <= n6223;
   BU20456_I(14) <= n6224;
   BU20456_I(15) <= n6225;
   BU20456_I(16) <= n6226;
   BU20456_I(17) <= n6227;
   BU20456_I(18) <= n6228;
   BU20456_I(19) <= n6229;
   BU20456_I(20) <= n6230;
   BU20456_I(21) <= n6231;
   BU20456_I(22) <= n6232;
   BU20456_I(23) <= n6233;
   BU20456_I(24) <= n6234;
   BU20456_I(25) <= n6235;
   n6405 <= BU20456_O;
   BU20456 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 26,
         c_input_inv_mask => "01111111111111111111111111"
      )
      PORT MAP (
         I => BU20456_I,
         O => BU20456_O
      );

   BU20487_I0 <= n6236;
   BU20487_I1 <= n6235;
   BU20487_I2 <= n6405;
   BU20487_I3 <= '0';
   n6402 <= BU20487_O;
   BU20487 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU20487_I0,
         I1 => BU20487_I1,
         I2 => BU20487_I2,
         I3 => BU20487_I3,
         O => BU20487_O
      );

   BU20488_A(0) <= n6236;
   BU20488_A(1) <= n6237;
   BU20488_A(2) <= n6238;
   BU20488_A(3) <= n6239;
   BU20488_A(4) <= n6240;
   BU20488_A(5) <= n6241;
   BU20488_A(6) <= n6242;
   BU20488_A(7) <= n6243;
   BU20488_A(8) <= n6244;
   BU20488_A(9) <= n6245;
   BU20488_A(10) <= n6246;
   BU20488_A(11) <= n6247;
   BU20488_A(12) <= n6248;
   BU20488_A(13) <= n6249;
   BU20488_A(14) <= n6250;
   BU20488_A(15) <= n6251;
   BU20488_B(0) <= n6402;
   n6385 <= BU20488_S(0);
   n6386 <= BU20488_S(1);
   n6387 <= BU20488_S(2);
   n6388 <= BU20488_S(3);
   n6389 <= BU20488_S(4);
   n6390 <= BU20488_S(5);
   n6391 <= BU20488_S(6);
   n6392 <= BU20488_S(7);
   n6393 <= BU20488_S(8);
   n6394 <= BU20488_S(9);
   n6395 <= BU20488_S(10);
   n6396 <= BU20488_S(11);
   n6397 <= BU20488_S(12);
   n6398 <= BU20488_S(13);
   n6399 <= BU20488_S(14);
   n6400 <= BU20488_S(15);
   BU20488 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 16,
         c_latency => 1,
         c_sinit_val => "00000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "00000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 17,
         c_low_bit => 0,
         c_ainit_val => "00000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 16,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU20488_A,
         B => BU20488_B,
         S => BU20488_S
      );

   BU20557_I0 <= n6251;
   BU20557_I1 <= n6250;
   BU20557_I2 <= n6400;
   BU20557_I3 <= '0';
   n6432 <= BU20557_O;
   BU20557 : LUT4
      GENERIC MAP (
         INIT  => X"0202"
      )
      PORT MAP (
         I0 => BU20557_I0,
         I1 => BU20557_I1,
         I2 => BU20557_I2,
         I3 => BU20557_I3,
         O => BU20557_O
      );

   BU20559_I0 <= n6251;
   BU20559_I1 <= n6400;
   BU20559_I2 <= '0';
   BU20559_I3 <= '0';
   n6434 <= BU20559_O;
   BU20559 : LUT4
      GENERIC MAP (
         INIT  => X"4444"
      )
      PORT MAP (
         I0 => BU20559_I0,
         I1 => BU20559_I1,
         I2 => BU20559_I2,
         I3 => BU20559_I3,
         O => BU20559_O
      );

   BU20560_D(0) <= n6385;
   BU20560_D(1) <= n6386;
   BU20560_D(2) <= n6387;
   BU20560_D(3) <= n6388;
   BU20560_D(4) <= n6389;
   BU20560_D(5) <= n6390;
   BU20560_D(6) <= n6391;
   BU20560_D(7) <= n6392;
   BU20560_D(8) <= n6393;
   BU20560_D(9) <= n6394;
   BU20560_D(10) <= n6395;
   BU20560_D(11) <= n6396;
   BU20560_D(12) <= n6397;
   BU20560_D(13) <= n6398;
   BU20560_D(14) <= n6399;
   n80 <= BU20560_Q(0);
   n81 <= BU20560_Q(1);
   n82 <= BU20560_Q(2);
   n83 <= BU20560_Q(3);
   n84 <= BU20560_Q(4);
   n85 <= BU20560_Q(5);
   n86 <= BU20560_Q(6);
   n87 <= BU20560_Q(7);
   n88 <= BU20560_Q(8);
   n89 <= BU20560_Q(9);
   n90 <= BU20560_Q(10);
   n91 <= BU20560_Q(11);
   n92 <= BU20560_Q(12);
   n93 <= BU20560_Q(13);
   n94 <= BU20560_Q(14);
   BU20560_CLK <= n152;
   BU20560_SCLR <= n6432;
   BU20560_SSET <= n6434;
   BU20560 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 15,
         c_has_ce => 0,
         c_sinit_val => "000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU20560_D,
         Q => BU20560_Q,
         CLK => BU20560_CLK,
         SCLR => BU20560_SCLR,
         SSET => BU20560_SSET
      );

   BU20621_D(0) <= n6400;
   n95 <= BU20621_Q(0);
   BU20621_CLK <= n152;
   BU20621_SCLR <= n6434;
   BU20621_SSET <= n6432;
   BU20621 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 0,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU20621_D,
         Q => BU20621_Q,
         CLK => BU20621_CLK,
         SCLR => BU20621_SCLR,
         SSET => BU20621_SSET
      );

   BU20628_D <= n6252;
   BU20628_C <= n152;
   BU20628_CE <= '1';
   n96 <= BU20628_Q;
   BU20628 : FDE
      PORT MAP (
         D => BU20628_D,
         C => BU20628_C,
         CE => BU20628_CE,
         Q => BU20628_Q
      );

   BU20631_ND <= n96;
   n131 <= BU20631_RDY;
   BU20631_CLK <= n152;
   BU20631_DIN(0) <= n80;
   BU20631_DIN(1) <= n81;
   BU20631_DIN(2) <= n82;
   BU20631_DIN(3) <= n83;
   BU20631_DIN(4) <= n84;
   BU20631_DIN(5) <= n85;
   BU20631_DIN(6) <= n86;
   BU20631_DIN(7) <= n87;
   BU20631_DIN(8) <= n88;
   BU20631_DIN(9) <= n89;
   BU20631_DIN(10) <= n90;
   BU20631_DIN(11) <= n91;
   BU20631_DIN(12) <= n92;
   BU20631_DIN(13) <= n93;
   BU20631_DIN(14) <= n94;
   BU20631_DIN(15) <= n95;
   n132 <= BU20631_SEL_O(0);
   n97 <= BU20631_DOUT(0);
   n98 <= BU20631_DOUT(1);
   n99 <= BU20631_DOUT(2);
   n100 <= BU20631_DOUT(3);
   n101 <= BU20631_DOUT(4);
   n102 <= BU20631_DOUT(5);
   n103 <= BU20631_DOUT(6);
   n104 <= BU20631_DOUT(7);
   n105 <= BU20631_DOUT(8);
   n106 <= BU20631_DOUT(9);
   n107 <= BU20631_DOUT(10);
   n108 <= BU20631_DOUT(11);
   n109 <= BU20631_DOUT(12);
   n110 <= BU20631_DOUT(13);
   n111 <= BU20631_DOUT(14);
   n112 <= BU20631_DOUT(15);
   n113 <= BU20631_DOUT(16);
   n114 <= BU20631_DOUT(17);
   n115 <= BU20631_DOUT(18);
   n116 <= BU20631_DOUT(19);
   n117 <= BU20631_DOUT(20);
   n118 <= BU20631_DOUT(21);
   n119 <= BU20631_DOUT(22);
   n120 <= BU20631_DOUT(23);
   n121 <= BU20631_DOUT(24);
   n122 <= BU20631_DOUT(25);
   n123 <= BU20631_DOUT(26);
   n124 <= BU20631_DOUT(27);
   n125 <= BU20631_DOUT(28);
   n126 <= BU20631_DOUT(29);
   n127 <= BU20631_DOUT(30);
   n128 <= BU20631_DOUT(31);
   n129 <= BU20631_DOUT(32);
   n130 <= BU20631_DOUT(33);
   BU20631 : C_DA_FIR_V7_0
      GENERIC MAP (
         c_has_sout_r => 0,
         c_result_width => 34,
         c_reload_delay => 657,
         c_data_type => 0,
         c_filter_type => 2,
         c_channels => 2,
         c_response => 0,
         c_has_sout_f => 0,
         c_reg_output => 0,
         c_taps => 66,
         c_data_width => 16,
         c_enable_rlocs => 0,
         c_coeff_type => 0,
         c_reload_mem_type => 2,
         c_has_sin_r => 0,
         c_reload => 0,
         c_baat => 1,
         c_latency => 26,
         c_coeff_width => 16,
         c_optimize => 1,
         c_use_model_func => 0,
         c_zpf => 1,
         c_has_sin_f => 0,
         c_shape => 0,
         c_saturate => 0,
         c_has_sel_o => 1,
         c_mem_init_file => "ddcv1_0_PFIR.mif",
         c_polyphase_factor => 5,
         c_has_sel_i => 0,
         c_has_reset => 0
      )
      PORT MAP (
         ND => BU20631_ND,
         RDY => BU20631_RDY,
         CLK => BU20631_CLK,
         RFD => BU20631_RFD,
         DIN => BU20631_DIN,
         SEL_O => BU20631_SEL_O,
         DOUT => BU20631_DOUT
      );

   BU24197_I0 <= n131;
   BU24197_I1 <= n132;
   BU24197_I2 <= '0';
   BU24197_I3 <= '0';
   n133 <= BU24197_O;
   BU24197 : LUT4
      GENERIC MAP (
         INIT  => X"2222"
      )
      PORT MAP (
         I0 => BU24197_I0,
         I1 => BU24197_I1,
         I2 => BU24197_I2,
         I3 => BU24197_I3,
         O => BU24197_O
      );

   BU24199_I0 <= n131;
   BU24199_I1 <= n132;
   BU24199_I2 <= '0';
   BU24199_I3 <= '0';
   n134 <= BU24199_O;
   BU24199 : LUT4
      GENERIC MAP (
         INIT  => X"8888"
      )
      PORT MAP (
         I0 => BU24199_I0,
         I1 => BU24199_I1,
         I2 => BU24199_I2,
         I3 => BU24199_I3,
         O => BU24199_O
      );

   BU24202_D <= n134;
   BU24202_C <= n152;
   BU24202_CE <= '1';
   n150 <= BU24202_Q;
   BU24202 : FDE
      PORT MAP (
         D => BU24202_D,
         C => BU24202_C,
         CE => BU24202_CE,
         Q => BU24202_Q
      );

   BU24207_I(0) <= n97;
   BU24207_I(1) <= n98;
   BU24207_I(2) <= n99;
   BU24207_I(3) <= n100;
   n6970 <= BU24207_O;
   BU24207 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 4,
         c_input_inv_mask => "0111"
      )
      PORT MAP (
         I => BU24207_I,
         O => BU24207_O
      );

   BU24213_I0 <= n101;
   BU24213_I1 <= n100;
   BU24213_I2 <= n6970;
   BU24213_I3 <= '0';
   n6967 <= BU24213_O;
   BU24213 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU24213_I0,
         I1 => BU24213_I1,
         I2 => BU24213_I2,
         I3 => BU24213_I3,
         O => BU24213_O
      );

   BU24214_A(0) <= n101;
   BU24214_A(1) <= n102;
   BU24214_A(2) <= n103;
   BU24214_A(3) <= n104;
   BU24214_A(4) <= n105;
   BU24214_A(5) <= n106;
   BU24214_A(6) <= n107;
   BU24214_A(7) <= n108;
   BU24214_A(8) <= n109;
   BU24214_A(9) <= n110;
   BU24214_A(10) <= n111;
   BU24214_A(11) <= n112;
   BU24214_A(12) <= n113;
   BU24214_A(13) <= n114;
   BU24214_A(14) <= n115;
   BU24214_A(15) <= n116;
   BU24214_A(16) <= n117;
   BU24214_A(17) <= n118;
   BU24214_A(18) <= n119;
   BU24214_A(19) <= n120;
   BU24214_A(20) <= n121;
   BU24214_A(21) <= n122;
   BU24214_A(22) <= n123;
   BU24214_A(23) <= n124;
   BU24214_A(24) <= n125;
   BU24214_A(25) <= n126;
   BU24214_A(26) <= n127;
   BU24214_A(27) <= n128;
   BU24214_A(28) <= n129;
   BU24214_A(29) <= n130;
   BU24214_B(0) <= n6967;
   n6936 <= BU24214_S(0);
   n6937 <= BU24214_S(1);
   n6938 <= BU24214_S(2);
   n6939 <= BU24214_S(3);
   n6940 <= BU24214_S(4);
   n6941 <= BU24214_S(5);
   n6942 <= BU24214_S(6);
   n6943 <= BU24214_S(7);
   n6944 <= BU24214_S(8);
   n6945 <= BU24214_S(9);
   n6946 <= BU24214_S(10);
   n6947 <= BU24214_S(11);
   n6948 <= BU24214_S(12);
   n6949 <= BU24214_S(13);
   n6950 <= BU24214_S(14);
   n6951 <= BU24214_S(15);
   n6952 <= BU24214_S(16);
   n6953 <= BU24214_S(17);
   n6954 <= BU24214_S(18);
   n6955 <= BU24214_S(19);
   n6956 <= BU24214_S(20);
   n6957 <= BU24214_S(21);
   n6958 <= BU24214_S(22);
   n6959 <= BU24214_S(23);
   n6960 <= BU24214_S(24);
   n6961 <= BU24214_S(25);
   n6962 <= BU24214_S(26);
   n6963 <= BU24214_S(27);
   n6964 <= BU24214_S(28);
   n6965 <= BU24214_S(29);
   BU24214 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 30,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 31,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 30,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU24214_A,
         B => BU24214_B,
         S => BU24214_S
      );

   BU24339_I0 <= n130;
   BU24339_I1 <= n129;
   BU24339_I2 <= n6965;
   BU24339_I3 <= n133;
   n6975 <= BU24339_O;
   BU24339 : LUT4
      GENERIC MAP (
         INIT  => X"0200"
      )
      PORT MAP (
         I0 => BU24339_I0,
         I1 => BU24339_I1,
         I2 => BU24339_I2,
         I3 => BU24339_I3,
         O => BU24339_O
      );

   BU24341_I0 <= n130;
   BU24341_I1 <= n6965;
   BU24341_I2 <= n133;
   BU24341_I3 <= '0';
   n6977 <= BU24341_O;
   BU24341 : LUT4
      GENERIC MAP (
         INIT  => X"4040"
      )
      PORT MAP (
         I0 => BU24341_I0,
         I1 => BU24341_I1,
         I2 => BU24341_I2,
         I3 => BU24341_I3,
         O => BU24341_O
      );

   BU24342_D(0) <= n6936;
   BU24342_D(1) <= n6937;
   BU24342_D(2) <= n6938;
   BU24342_D(3) <= n6939;
   BU24342_D(4) <= n6940;
   BU24342_D(5) <= n6941;
   BU24342_D(6) <= n6942;
   BU24342_D(7) <= n6943;
   BU24342_D(8) <= n6944;
   BU24342_D(9) <= n6945;
   BU24342_D(10) <= n6946;
   BU24342_D(11) <= n6947;
   BU24342_D(12) <= n6948;
   BU24342_D(13) <= n6949;
   BU24342_D(14) <= n6950;
   BU24342_D(15) <= n6951;
   BU24342_D(16) <= n6952;
   BU24342_D(17) <= n6953;
   BU24342_D(18) <= n6954;
   BU24342_D(19) <= n6955;
   BU24342_D(20) <= n6956;
   BU24342_D(21) <= n6957;
   BU24342_D(22) <= n6958;
   BU24342_D(23) <= n6959;
   BU24342_D(24) <= n6960;
   BU24342_D(25) <= n6961;
   BU24342_D(26) <= n6962;
   BU24342_D(27) <= n6963;
   BU24342_D(28) <= n6964;
   n192 <= BU24342_Q(0);
   n193 <= BU24342_Q(1);
   n194 <= BU24342_Q(2);
   n195 <= BU24342_Q(3);
   n196 <= BU24342_Q(4);
   n197 <= BU24342_Q(5);
   n198 <= BU24342_Q(6);
   n199 <= BU24342_Q(7);
   n200 <= BU24342_Q(8);
   n201 <= BU24342_Q(9);
   n202 <= BU24342_Q(10);
   n203 <= BU24342_Q(11);
   n204 <= BU24342_Q(12);
   n205 <= BU24342_Q(13);
   n206 <= BU24342_Q(14);
   n207 <= BU24342_Q(15);
   n208 <= BU24342_Q(16);
   n209 <= BU24342_Q(17);
   n210 <= BU24342_Q(18);
   n211 <= BU24342_Q(19);
   n212 <= BU24342_Q(20);
   n213 <= BU24342_Q(21);
   n214 <= BU24342_Q(22);
   n215 <= BU24342_Q(23);
   n216 <= BU24342_Q(24);
   n217 <= BU24342_Q(25);
   n218 <= BU24342_Q(26);
   n219 <= BU24342_Q(27);
   n220 <= BU24342_Q(28);
   BU24342_CLK <= n152;
   BU24342_CE <= n133;
   BU24342_SCLR <= n6975;
   BU24342_SSET <= n6977;
   BU24342 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 29,
         c_has_ce => 1,
         c_sinit_val => "00000000000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU24342_D,
         Q => BU24342_Q,
         CLK => BU24342_CLK,
         CE => BU24342_CE,
         SCLR => BU24342_SCLR,
         SSET => BU24342_SSET
      );

   BU24462_D(0) <= n6965;
   n221 <= BU24462_Q(0);
   BU24462_CLK <= n152;
   BU24462_CE <= n133;
   BU24462_SCLR <= n6977;
   BU24462_SSET <= n6975;
   BU24462 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 1,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU24462_D,
         Q => BU24462_Q,
         CLK => BU24462_CLK,
         CE => BU24462_CE,
         SCLR => BU24462_SCLR,
         SSET => BU24462_SSET
      );

   BU24474_I(0) <= n97;
   BU24474_I(1) <= n98;
   BU24474_I(2) <= n99;
   BU24474_I(3) <= n100;
   n7511 <= BU24474_O;
   BU24474 : C_GATE_BIT_V5_0
      GENERIC MAP (
         c_has_aset => 0,
         c_gate_type => 0,
         c_sync_priority => 1,
         c_has_sclr => 0,
         c_enable_rlocs => 0,
         c_ainit_val => "0",
         c_pipe_stages => 0,
         c_has_ce => 0,
         c_has_aclr => 0,
         c_sync_enable => 0,
         c_has_ainit => 0,
         c_sinit_val => "0",
         c_has_sset => 0,
         c_has_sinit => 0,
         c_has_q => 0,
         c_has_o => 1,
         c_inputs => 4,
         c_input_inv_mask => "0111"
      )
      PORT MAP (
         I => BU24474_I,
         O => BU24474_O
      );

   BU24480_I0 <= n101;
   BU24480_I1 <= n100;
   BU24480_I2 <= n7511;
   BU24480_I3 <= '0';
   n7508 <= BU24480_O;
   BU24480 : LUT4
      GENERIC MAP (
         INIT  => X"8c8c"
      )
      PORT MAP (
         I0 => BU24480_I0,
         I1 => BU24480_I1,
         I2 => BU24480_I2,
         I3 => BU24480_I3,
         O => BU24480_O
      );

   BU24481_A(0) <= n101;
   BU24481_A(1) <= n102;
   BU24481_A(2) <= n103;
   BU24481_A(3) <= n104;
   BU24481_A(4) <= n105;
   BU24481_A(5) <= n106;
   BU24481_A(6) <= n107;
   BU24481_A(7) <= n108;
   BU24481_A(8) <= n109;
   BU24481_A(9) <= n110;
   BU24481_A(10) <= n111;
   BU24481_A(11) <= n112;
   BU24481_A(12) <= n113;
   BU24481_A(13) <= n114;
   BU24481_A(14) <= n115;
   BU24481_A(15) <= n116;
   BU24481_A(16) <= n117;
   BU24481_A(17) <= n118;
   BU24481_A(18) <= n119;
   BU24481_A(19) <= n120;
   BU24481_A(20) <= n121;
   BU24481_A(21) <= n122;
   BU24481_A(22) <= n123;
   BU24481_A(23) <= n124;
   BU24481_A(24) <= n125;
   BU24481_A(25) <= n126;
   BU24481_A(26) <= n127;
   BU24481_A(27) <= n128;
   BU24481_A(28) <= n129;
   BU24481_A(29) <= n130;
   BU24481_B(0) <= n7508;
   n7477 <= BU24481_S(0);
   n7478 <= BU24481_S(1);
   n7479 <= BU24481_S(2);
   n7480 <= BU24481_S(3);
   n7481 <= BU24481_S(4);
   n7482 <= BU24481_S(5);
   n7483 <= BU24481_S(6);
   n7484 <= BU24481_S(7);
   n7485 <= BU24481_S(8);
   n7486 <= BU24481_S(9);
   n7487 <= BU24481_S(10);
   n7488 <= BU24481_S(11);
   n7489 <= BU24481_S(12);
   n7490 <= BU24481_S(13);
   n7491 <= BU24481_S(14);
   n7492 <= BU24481_S(15);
   n7493 <= BU24481_S(16);
   n7494 <= BU24481_S(17);
   n7495 <= BU24481_S(18);
   n7496 <= BU24481_S(19);
   n7497 <= BU24481_S(20);
   n7498 <= BU24481_S(21);
   n7499 <= BU24481_S(22);
   n7500 <= BU24481_S(23);
   n7501 <= BU24481_S(24);
   n7502 <= BU24481_S(25);
   n7503 <= BU24481_S(26);
   n7504 <= BU24481_S(27);
   n7505 <= BU24481_S(28);
   n7506 <= BU24481_S(29);
   BU24481 : C_ADDSUB_V5_0
      GENERIC MAP (
         c_has_bypass_with_cin => 0,
         c_a_type => 0,
         c_has_sclr => 0,
         c_has_aset => 0,
         c_has_b_out => 0,
         c_sync_priority => 1,
         c_has_s => 1,
         c_has_q => 0,
         c_bypass_enable => 0,
         c_b_constant => 0,
         c_has_ovfl => 0,
         c_high_bit => 30,
         c_latency => 1,
         c_sinit_val => "0000000000000000000000000000000",
         c_has_bypass => 0,
         c_pipe_stages => 0,
         c_has_sset => 0,
         c_has_ainit => 0,
         c_has_a_signed => 0,
         c_has_q_c_out => 0,
         c_b_type => 1,
         c_has_add => 0,
         c_has_sinit => 0,
         c_has_b_in => 0,
         c_has_b_signed => 0,
         c_bypass_low => 0,
         c_enable_rlocs => 0,
         c_b_value => "0000000000000000000000000000000",
         c_add_mode => 0,
         c_has_aclr => 0,
         c_out_width => 31,
         c_low_bit => 0,
         c_ainit_val => "0000000000000000000000000000000",
         c_has_q_ovfl => 0,
         c_has_q_b_out => 0,
         c_has_c_out => 0,
         c_b_width => 1,
         c_a_width => 30,
         c_sync_enable => 0,
         c_has_ce => 0,
         c_has_c_in => 0
      )
      PORT MAP (
         A => BU24481_A,
         B => BU24481_B,
         S => BU24481_S
      );

   BU24606_I0 <= n130;
   BU24606_I1 <= n129;
   BU24606_I2 <= n7506;
   BU24606_I3 <= n134;
   n7516 <= BU24606_O;
   BU24606 : LUT4
      GENERIC MAP (
         INIT  => X"0200"
      )
      PORT MAP (
         I0 => BU24606_I0,
         I1 => BU24606_I1,
         I2 => BU24606_I2,
         I3 => BU24606_I3,
         O => BU24606_O
      );

   BU24608_I0 <= n130;
   BU24608_I1 <= n7506;
   BU24608_I2 <= n134;
   BU24608_I3 <= '0';
   n7518 <= BU24608_O;
   BU24608 : LUT4
      GENERIC MAP (
         INIT  => X"4040"
      )
      PORT MAP (
         I0 => BU24608_I0,
         I1 => BU24608_I1,
         I2 => BU24608_I2,
         I3 => BU24608_I3,
         O => BU24608_O
      );

   BU24609_D(0) <= n7477;
   BU24609_D(1) <= n7478;
   BU24609_D(2) <= n7479;
   BU24609_D(3) <= n7480;
   BU24609_D(4) <= n7481;
   BU24609_D(5) <= n7482;
   BU24609_D(6) <= n7483;
   BU24609_D(7) <= n7484;
   BU24609_D(8) <= n7485;
   BU24609_D(9) <= n7486;
   BU24609_D(10) <= n7487;
   BU24609_D(11) <= n7488;
   BU24609_D(12) <= n7489;
   BU24609_D(13) <= n7490;
   BU24609_D(14) <= n7491;
   BU24609_D(15) <= n7492;
   BU24609_D(16) <= n7493;
   BU24609_D(17) <= n7494;
   BU24609_D(18) <= n7495;
   BU24609_D(19) <= n7496;
   BU24609_D(20) <= n7497;
   BU24609_D(21) <= n7498;
   BU24609_D(22) <= n7499;
   BU24609_D(23) <= n7500;
   BU24609_D(24) <= n7501;
   BU24609_D(25) <= n7502;
   BU24609_D(26) <= n7503;
   BU24609_D(27) <= n7504;
   BU24609_D(28) <= n7505;
   n222 <= BU24609_Q(0);
   n223 <= BU24609_Q(1);
   n224 <= BU24609_Q(2);
   n225 <= BU24609_Q(3);
   n226 <= BU24609_Q(4);
   n227 <= BU24609_Q(5);
   n228 <= BU24609_Q(6);
   n229 <= BU24609_Q(7);
   n230 <= BU24609_Q(8);
   n231 <= BU24609_Q(9);
   n232 <= BU24609_Q(10);
   n233 <= BU24609_Q(11);
   n234 <= BU24609_Q(12);
   n235 <= BU24609_Q(13);
   n236 <= BU24609_Q(14);
   n237 <= BU24609_Q(15);
   n238 <= BU24609_Q(16);
   n239 <= BU24609_Q(17);
   n240 <= BU24609_Q(18);
   n241 <= BU24609_Q(19);
   n242 <= BU24609_Q(20);
   n243 <= BU24609_Q(21);
   n244 <= BU24609_Q(22);
   n245 <= BU24609_Q(23);
   n246 <= BU24609_Q(24);
   n247 <= BU24609_Q(25);
   n248 <= BU24609_Q(26);
   n249 <= BU24609_Q(27);
   n250 <= BU24609_Q(28);
   BU24609_CLK <= n152;
   BU24609_CE <= n134;
   BU24609_SCLR <= n7516;
   BU24609_SSET <= n7518;
   BU24609 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 29,
         c_has_ce => 1,
         c_sinit_val => "00000000000000000000000000000",
         c_has_sinit => 0,
         c_ainit_val => "00000000000000000000000000000",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU24609_D,
         Q => BU24609_Q,
         CLK => BU24609_CLK,
         CE => BU24609_CE,
         SCLR => BU24609_SCLR,
         SSET => BU24609_SSET
      );

   BU24729_D(0) <= n7506;
   n251 <= BU24729_Q(0);
   BU24729_CLK <= n152;
   BU24729_CE <= n134;
   BU24729_SCLR <= n7518;
   BU24729_SSET <= n7516;
   BU24729 : C_REG_FD_V5_0
      GENERIC MAP (
         c_width => 1,
         c_has_ce => 1,
         c_sinit_val => "0",
         c_has_sinit => 0,
         c_ainit_val => "0",
         c_has_aset => 0,
         c_sync_enable => 0,
         c_enable_rlocs => 0,
         c_has_aclr => 0,
         c_has_sset => 1,
         c_sync_priority => 0,
         c_has_ainit => 0,
         c_has_sclr => 1
      )
      PORT MAP (
         D => BU24729_D,
         Q => BU24729_Q,
         CLK => BU24729_CLK,
         CE => BU24729_CE,
         SCLR => BU24729_SCLR,
         SSET => BU24729_SSET
      );


END xilinx;


-- synopsys translate_on
